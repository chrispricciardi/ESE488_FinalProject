
module sigmoid ( clk, reset, done, d, we, sig_ready, sig_in, address, sig_out
 );
  input [15:0] d;
  input [15:0] sig_in;
  input [6:0] address;
  output [15:0] sig_out;
  input clk, reset, done, we;
  output sig_ready;
  wire   \x[120][15] , \x[120][14] , \x[120][13] , \x[120][12] , \x[120][11] ,
         \x[120][10] , \x[120][9] , \x[120][8] , \x[120][7] , \x[120][6] ,
         \x[120][5] , \x[120][4] , \x[120][3] , \x[120][2] , \x[120][1] ,
         \x[120][0] , \x[119][15] , \x[119][14] , \x[119][13] , \x[119][12] ,
         \x[119][11] , \x[119][10] , \x[119][9] , \x[119][8] , \x[119][7] ,
         \x[119][6] , \x[119][5] , \x[119][4] , \x[119][3] , \x[119][2] ,
         \x[119][1] , \x[119][0] , \x[118][15] , \x[118][14] , \x[118][13] ,
         \x[118][12] , \x[118][11] , \x[118][10] , \x[118][9] , \x[118][8] ,
         \x[118][7] , \x[118][6] , \x[118][5] , \x[118][4] , \x[118][3] ,
         \x[118][2] , \x[118][1] , \x[118][0] , \x[117][15] , \x[117][14] ,
         \x[117][13] , \x[117][12] , \x[117][11] , \x[117][10] , \x[117][9] ,
         \x[117][8] , \x[117][7] , \x[117][6] , \x[117][5] , \x[117][4] ,
         \x[117][3] , \x[117][2] , \x[117][1] , \x[117][0] , \x[116][15] ,
         \x[116][14] , \x[116][13] , \x[116][12] , \x[116][11] , \x[116][10] ,
         \x[116][9] , \x[116][8] , \x[116][7] , \x[116][6] , \x[116][5] ,
         \x[116][4] , \x[116][3] , \x[116][2] , \x[116][1] , \x[116][0] ,
         \x[115][15] , \x[115][14] , \x[115][13] , \x[115][12] , \x[115][11] ,
         \x[115][10] , \x[115][9] , \x[115][8] , \x[115][7] , \x[115][6] ,
         \x[115][5] , \x[115][4] , \x[115][3] , \x[115][2] , \x[115][1] ,
         \x[115][0] , \x[114][15] , \x[114][14] , \x[114][13] , \x[114][12] ,
         \x[114][11] , \x[114][10] , \x[114][9] , \x[114][8] , \x[114][7] ,
         \x[114][6] , \x[114][5] , \x[114][4] , \x[114][3] , \x[114][2] ,
         \x[114][1] , \x[114][0] , \x[113][15] , \x[113][14] , \x[113][13] ,
         \x[113][12] , \x[113][11] , \x[113][10] , \x[113][9] , \x[113][8] ,
         \x[113][7] , \x[113][6] , \x[113][5] , \x[113][4] , \x[113][3] ,
         \x[113][2] , \x[113][1] , \x[113][0] , \x[112][15] , \x[112][14] ,
         \x[112][13] , \x[112][12] , \x[112][11] , \x[112][10] , \x[112][9] ,
         \x[112][8] , \x[112][7] , \x[112][6] , \x[112][5] , \x[112][4] ,
         \x[112][3] , \x[112][2] , \x[112][1] , \x[112][0] , \x[111][15] ,
         \x[111][14] , \x[111][13] , \x[111][12] , \x[111][11] , \x[111][10] ,
         \x[111][9] , \x[111][8] , \x[111][7] , \x[111][6] , \x[111][5] ,
         \x[111][4] , \x[111][3] , \x[111][2] , \x[111][1] , \x[111][0] ,
         \x[110][15] , \x[110][14] , \x[110][13] , \x[110][12] , \x[110][11] ,
         \x[110][10] , \x[110][9] , \x[110][8] , \x[110][7] , \x[110][6] ,
         \x[110][5] , \x[110][4] , \x[110][3] , \x[110][2] , \x[110][1] ,
         \x[110][0] , \x[109][15] , \x[109][14] , \x[109][13] , \x[109][12] ,
         \x[109][11] , \x[109][10] , \x[109][9] , \x[109][8] , \x[109][7] ,
         \x[109][6] , \x[109][5] , \x[109][4] , \x[109][3] , \x[109][2] ,
         \x[109][1] , \x[109][0] , \x[108][15] , \x[108][14] , \x[108][13] ,
         \x[108][12] , \x[108][11] , \x[108][10] , \x[108][9] , \x[108][8] ,
         \x[108][7] , \x[108][6] , \x[108][5] , \x[108][4] , \x[108][3] ,
         \x[108][2] , \x[108][1] , \x[108][0] , \x[107][15] , \x[107][14] ,
         \x[107][13] , \x[107][12] , \x[107][11] , \x[107][10] , \x[107][9] ,
         \x[107][8] , \x[107][7] , \x[107][6] , \x[107][5] , \x[107][4] ,
         \x[107][3] , \x[107][2] , \x[107][1] , \x[107][0] , \x[106][15] ,
         \x[106][14] , \x[106][13] , \x[106][12] , \x[106][11] , \x[106][10] ,
         \x[106][9] , \x[106][8] , \x[106][7] , \x[106][6] , \x[106][5] ,
         \x[106][4] , \x[106][3] , \x[106][2] , \x[106][1] , \x[106][0] ,
         \x[105][15] , \x[105][14] , \x[105][13] , \x[105][12] , \x[105][11] ,
         \x[105][10] , \x[105][9] , \x[105][8] , \x[105][7] , \x[105][6] ,
         \x[105][5] , \x[105][4] , \x[105][3] , \x[105][2] , \x[105][1] ,
         \x[105][0] , \x[104][15] , \x[104][14] , \x[104][13] , \x[104][12] ,
         \x[104][11] , \x[104][10] , \x[104][9] , \x[104][8] , \x[104][7] ,
         \x[104][6] , \x[104][5] , \x[104][4] , \x[104][3] , \x[104][2] ,
         \x[104][1] , \x[104][0] , \x[103][15] , \x[103][14] , \x[103][13] ,
         \x[103][12] , \x[103][11] , \x[103][10] , \x[103][9] , \x[103][8] ,
         \x[103][7] , \x[103][6] , \x[103][5] , \x[103][4] , \x[103][3] ,
         \x[103][2] , \x[103][1] , \x[103][0] , \x[102][15] , \x[102][14] ,
         \x[102][13] , \x[102][12] , \x[102][11] , \x[102][10] , \x[102][9] ,
         \x[102][8] , \x[102][7] , \x[102][6] , \x[102][5] , \x[102][4] ,
         \x[102][3] , \x[102][2] , \x[102][1] , \x[102][0] , \x[101][15] ,
         \x[101][14] , \x[101][13] , \x[101][12] , \x[101][11] , \x[101][10] ,
         \x[101][9] , \x[101][8] , \x[101][7] , \x[101][6] , \x[101][5] ,
         \x[101][4] , \x[101][3] , \x[101][2] , \x[101][1] , \x[101][0] ,
         \x[100][15] , \x[100][14] , \x[100][13] , \x[100][12] , \x[100][11] ,
         \x[100][10] , \x[100][9] , \x[100][8] , \x[100][7] , \x[100][6] ,
         \x[100][5] , \x[100][4] , \x[100][3] , \x[100][2] , \x[100][1] ,
         \x[100][0] , \x[99][15] , \x[99][14] , \x[99][13] , \x[99][12] ,
         \x[99][11] , \x[99][10] , \x[99][9] , \x[99][8] , \x[99][7] ,
         \x[99][6] , \x[99][5] , \x[99][4] , \x[99][3] , \x[99][2] ,
         \x[99][1] , \x[99][0] , \x[98][15] , \x[98][14] , \x[98][13] ,
         \x[98][12] , \x[98][11] , \x[98][10] , \x[98][9] , \x[98][8] ,
         \x[98][7] , \x[98][6] , \x[98][5] , \x[98][4] , \x[98][3] ,
         \x[98][2] , \x[98][1] , \x[98][0] , \x[97][15] , \x[97][14] ,
         \x[97][13] , \x[97][12] , \x[97][11] , \x[97][10] , \x[97][9] ,
         \x[97][8] , \x[97][7] , \x[97][6] , \x[97][5] , \x[97][4] ,
         \x[97][3] , \x[97][2] , \x[97][1] , \x[97][0] , \x[96][15] ,
         \x[96][14] , \x[96][13] , \x[96][12] , \x[96][11] , \x[96][10] ,
         \x[96][9] , \x[96][8] , \x[96][7] , \x[96][6] , \x[96][5] ,
         \x[96][4] , \x[96][3] , \x[96][2] , \x[96][1] , \x[96][0] ,
         \x[95][15] , \x[95][14] , \x[95][13] , \x[95][12] , \x[95][11] ,
         \x[95][10] , \x[95][9] , \x[95][8] , \x[95][7] , \x[95][6] ,
         \x[95][5] , \x[95][4] , \x[95][3] , \x[95][2] , \x[95][1] ,
         \x[95][0] , \x[94][15] , \x[94][14] , \x[94][13] , \x[94][12] ,
         \x[94][11] , \x[94][10] , \x[94][9] , \x[94][8] , \x[94][7] ,
         \x[94][6] , \x[94][5] , \x[94][4] , \x[94][3] , \x[94][2] ,
         \x[94][1] , \x[94][0] , \x[93][15] , \x[93][14] , \x[93][13] ,
         \x[93][12] , \x[93][11] , \x[93][10] , \x[93][9] , \x[93][8] ,
         \x[93][7] , \x[93][6] , \x[93][5] , \x[93][4] , \x[93][3] ,
         \x[93][2] , \x[93][1] , \x[93][0] , \x[92][15] , \x[92][14] ,
         \x[92][13] , \x[92][12] , \x[92][11] , \x[92][10] , \x[92][9] ,
         \x[92][8] , \x[92][7] , \x[92][6] , \x[92][5] , \x[92][4] ,
         \x[92][3] , \x[92][2] , \x[92][1] , \x[92][0] , \x[91][15] ,
         \x[91][14] , \x[91][13] , \x[91][12] , \x[91][11] , \x[91][10] ,
         \x[91][9] , \x[91][8] , \x[91][7] , \x[91][6] , \x[91][5] ,
         \x[91][4] , \x[91][3] , \x[91][2] , \x[91][1] , \x[91][0] ,
         \x[90][15] , \x[90][14] , \x[90][13] , \x[90][12] , \x[90][11] ,
         \x[90][10] , \x[90][9] , \x[90][8] , \x[90][7] , \x[90][6] ,
         \x[90][5] , \x[90][4] , \x[90][3] , \x[90][2] , \x[90][1] ,
         \x[90][0] , \x[89][15] , \x[89][14] , \x[89][13] , \x[89][12] ,
         \x[89][11] , \x[89][10] , \x[89][9] , \x[89][8] , \x[89][7] ,
         \x[89][6] , \x[89][5] , \x[89][4] , \x[89][3] , \x[89][2] ,
         \x[89][1] , \x[89][0] , \x[88][15] , \x[88][14] , \x[88][13] ,
         \x[88][12] , \x[88][11] , \x[88][10] , \x[88][9] , \x[88][8] ,
         \x[88][7] , \x[88][6] , \x[88][5] , \x[88][4] , \x[88][3] ,
         \x[88][2] , \x[88][1] , \x[88][0] , \x[87][15] , \x[87][14] ,
         \x[87][13] , \x[87][12] , \x[87][11] , \x[87][10] , \x[87][9] ,
         \x[87][8] , \x[87][7] , \x[87][6] , \x[87][5] , \x[87][4] ,
         \x[87][3] , \x[87][2] , \x[87][1] , \x[87][0] , \x[86][15] ,
         \x[86][14] , \x[86][13] , \x[86][12] , \x[86][11] , \x[86][10] ,
         \x[86][9] , \x[86][8] , \x[86][7] , \x[86][6] , \x[86][5] ,
         \x[86][4] , \x[86][3] , \x[86][2] , \x[86][1] , \x[86][0] ,
         \x[85][15] , \x[85][14] , \x[85][13] , \x[85][12] , \x[85][11] ,
         \x[85][10] , \x[85][9] , \x[85][8] , \x[85][7] , \x[85][6] ,
         \x[85][5] , \x[85][4] , \x[85][3] , \x[85][2] , \x[85][1] ,
         \x[85][0] , \x[84][15] , \x[84][14] , \x[84][13] , \x[84][12] ,
         \x[84][11] , \x[84][10] , \x[84][9] , \x[84][8] , \x[84][7] ,
         \x[84][6] , \x[84][5] , \x[84][4] , \x[84][3] , \x[84][2] ,
         \x[84][1] , \x[84][0] , \x[83][15] , \x[83][14] , \x[83][13] ,
         \x[83][12] , \x[83][11] , \x[83][10] , \x[83][9] , \x[83][8] ,
         \x[83][7] , \x[83][6] , \x[83][5] , \x[83][4] , \x[83][3] ,
         \x[83][2] , \x[83][1] , \x[83][0] , \x[82][15] , \x[82][14] ,
         \x[82][13] , \x[82][12] , \x[82][11] , \x[82][10] , \x[82][9] ,
         \x[82][8] , \x[82][7] , \x[82][6] , \x[82][5] , \x[82][4] ,
         \x[82][3] , \x[82][2] , \x[82][1] , \x[82][0] , \x[81][15] ,
         \x[81][14] , \x[81][13] , \x[81][12] , \x[81][11] , \x[81][10] ,
         \x[81][9] , \x[81][8] , \x[81][7] , \x[81][6] , \x[81][5] ,
         \x[81][4] , \x[81][3] , \x[81][2] , \x[81][1] , \x[81][0] ,
         \x[80][15] , \x[80][14] , \x[80][13] , \x[80][12] , \x[80][11] ,
         \x[80][10] , \x[80][9] , \x[80][8] , \x[80][7] , \x[80][6] ,
         \x[80][5] , \x[80][4] , \x[80][3] , \x[80][2] , \x[80][1] ,
         \x[80][0] , \x[79][15] , \x[79][14] , \x[79][13] , \x[79][12] ,
         \x[79][11] , \x[79][10] , \x[79][9] , \x[79][8] , \x[79][7] ,
         \x[79][6] , \x[79][5] , \x[79][4] , \x[79][3] , \x[79][2] ,
         \x[79][1] , \x[79][0] , \x[78][15] , \x[78][14] , \x[78][13] ,
         \x[78][12] , \x[78][11] , \x[78][10] , \x[78][9] , \x[78][8] ,
         \x[78][7] , \x[78][6] , \x[78][5] , \x[78][4] , \x[78][3] ,
         \x[78][2] , \x[78][1] , \x[78][0] , \x[77][15] , \x[77][14] ,
         \x[77][13] , \x[77][12] , \x[77][11] , \x[77][10] , \x[77][9] ,
         \x[77][8] , \x[77][7] , \x[77][6] , \x[77][5] , \x[77][4] ,
         \x[77][3] , \x[77][2] , \x[77][1] , \x[77][0] , \x[76][15] ,
         \x[76][14] , \x[76][13] , \x[76][12] , \x[76][11] , \x[76][10] ,
         \x[76][9] , \x[76][8] , \x[76][7] , \x[76][6] , \x[76][5] ,
         \x[76][4] , \x[76][3] , \x[76][2] , \x[76][1] , \x[76][0] ,
         \x[75][15] , \x[75][14] , \x[75][13] , \x[75][12] , \x[75][11] ,
         \x[75][10] , \x[75][9] , \x[75][8] , \x[75][7] , \x[75][6] ,
         \x[75][5] , \x[75][4] , \x[75][3] , \x[75][2] , \x[75][1] ,
         \x[75][0] , \x[74][15] , \x[74][14] , \x[74][13] , \x[74][12] ,
         \x[74][11] , \x[74][10] , \x[74][9] , \x[74][8] , \x[74][7] ,
         \x[74][6] , \x[74][5] , \x[74][4] , \x[74][3] , \x[74][2] ,
         \x[74][1] , \x[74][0] , \x[73][15] , \x[73][14] , \x[73][13] ,
         \x[73][12] , \x[73][11] , \x[73][10] , \x[73][9] , \x[73][8] ,
         \x[73][7] , \x[73][6] , \x[73][5] , \x[73][4] , \x[73][3] ,
         \x[73][2] , \x[73][1] , \x[73][0] , \x[72][15] , \x[72][14] ,
         \x[72][13] , \x[72][12] , \x[72][11] , \x[72][10] , \x[72][9] ,
         \x[72][8] , \x[72][7] , \x[72][6] , \x[72][5] , \x[72][4] ,
         \x[72][3] , \x[72][2] , \x[72][1] , \x[72][0] , \x[71][15] ,
         \x[71][14] , \x[71][13] , \x[71][12] , \x[71][11] , \x[71][10] ,
         \x[71][9] , \x[71][8] , \x[71][7] , \x[71][6] , \x[71][5] ,
         \x[71][4] , \x[71][3] , \x[71][2] , \x[71][1] , \x[71][0] ,
         \x[70][15] , \x[70][14] , \x[70][13] , \x[70][12] , \x[70][11] ,
         \x[70][10] , \x[70][9] , \x[70][8] , \x[70][7] , \x[70][6] ,
         \x[70][5] , \x[70][4] , \x[70][3] , \x[70][2] , \x[70][1] ,
         \x[70][0] , \x[69][15] , \x[69][14] , \x[69][13] , \x[69][12] ,
         \x[69][11] , \x[69][10] , \x[69][9] , \x[69][8] , \x[69][7] ,
         \x[69][6] , \x[69][5] , \x[69][4] , \x[69][3] , \x[69][2] ,
         \x[69][1] , \x[69][0] , \x[68][15] , \x[68][14] , \x[68][13] ,
         \x[68][12] , \x[68][11] , \x[68][10] , \x[68][9] , \x[68][8] ,
         \x[68][7] , \x[68][6] , \x[68][5] , \x[68][4] , \x[68][3] ,
         \x[68][2] , \x[68][1] , \x[68][0] , \x[67][15] , \x[67][14] ,
         \x[67][13] , \x[67][12] , \x[67][11] , \x[67][10] , \x[67][9] ,
         \x[67][8] , \x[67][7] , \x[67][6] , \x[67][5] , \x[67][4] ,
         \x[67][3] , \x[67][2] , \x[67][1] , \x[67][0] , \x[66][15] ,
         \x[66][14] , \x[66][13] , \x[66][12] , \x[66][11] , \x[66][10] ,
         \x[66][9] , \x[66][8] , \x[66][7] , \x[66][6] , \x[66][5] ,
         \x[66][4] , \x[66][3] , \x[66][2] , \x[66][1] , \x[66][0] ,
         \x[65][15] , \x[65][14] , \x[65][13] , \x[65][12] , \x[65][11] ,
         \x[65][10] , \x[65][9] , \x[65][8] , \x[65][7] , \x[65][6] ,
         \x[65][5] , \x[65][4] , \x[65][3] , \x[65][2] , \x[65][1] ,
         \x[65][0] , \x[64][15] , \x[64][14] , \x[64][13] , \x[64][12] ,
         \x[64][11] , \x[64][10] , \x[64][9] , \x[64][8] , \x[64][7] ,
         \x[64][6] , \x[64][5] , \x[64][4] , \x[64][3] , \x[64][2] ,
         \x[64][1] , \x[64][0] , \x[63][15] , \x[63][14] , \x[63][13] ,
         \x[63][12] , \x[63][11] , \x[63][10] , \x[63][9] , \x[63][8] ,
         \x[63][7] , \x[63][6] , \x[63][5] , \x[63][4] , \x[63][3] ,
         \x[63][2] , \x[63][1] , \x[63][0] , \x[62][15] , \x[62][14] ,
         \x[62][13] , \x[62][12] , \x[62][11] , \x[62][10] , \x[62][9] ,
         \x[62][8] , \x[62][7] , \x[62][6] , \x[62][5] , \x[62][4] ,
         \x[62][3] , \x[62][2] , \x[62][1] , \x[62][0] , \x[61][15] ,
         \x[61][14] , \x[61][13] , \x[61][12] , \x[61][11] , \x[61][10] ,
         \x[61][9] , \x[61][8] , \x[61][7] , \x[61][6] , \x[61][5] ,
         \x[61][4] , \x[61][3] , \x[61][2] , \x[61][1] , \x[61][0] ,
         \x[60][15] , \x[60][14] , \x[60][13] , \x[60][12] , \x[60][11] ,
         \x[60][10] , \x[60][9] , \x[60][8] , \x[60][7] , \x[60][6] ,
         \x[60][5] , \x[60][4] , \x[60][3] , \x[60][2] , \x[60][1] ,
         \x[60][0] , \x[59][15] , \x[59][14] , \x[59][13] , \x[59][12] ,
         \x[59][11] , \x[59][10] , \x[59][9] , \x[59][8] , \x[59][7] ,
         \x[59][6] , \x[59][5] , \x[59][4] , \x[59][3] , \x[59][2] ,
         \x[59][1] , \x[59][0] , \x[58][15] , \x[58][14] , \x[58][13] ,
         \x[58][12] , \x[58][11] , \x[58][10] , \x[58][9] , \x[58][8] ,
         \x[58][7] , \x[58][6] , \x[58][5] , \x[58][4] , \x[58][3] ,
         \x[58][2] , \x[58][1] , \x[58][0] , \x[57][15] , \x[57][14] ,
         \x[57][13] , \x[57][12] , \x[57][11] , \x[57][10] , \x[57][9] ,
         \x[57][8] , \x[57][7] , \x[57][6] , \x[57][5] , \x[57][4] ,
         \x[57][3] , \x[57][2] , \x[57][1] , \x[57][0] , \x[56][15] ,
         \x[56][14] , \x[56][13] , \x[56][12] , \x[56][11] , \x[56][10] ,
         \x[56][9] , \x[56][8] , \x[56][7] , \x[56][6] , \x[56][5] ,
         \x[56][4] , \x[56][3] , \x[56][2] , \x[56][1] , \x[56][0] ,
         \x[55][15] , \x[55][14] , \x[55][13] , \x[55][12] , \x[55][11] ,
         \x[55][10] , \x[55][9] , \x[55][8] , \x[55][7] , \x[55][6] ,
         \x[55][5] , \x[55][4] , \x[55][3] , \x[55][2] , \x[55][1] ,
         \x[55][0] , \x[54][15] , \x[54][14] , \x[54][13] , \x[54][12] ,
         \x[54][11] , \x[54][10] , \x[54][9] , \x[54][8] , \x[54][7] ,
         \x[54][6] , \x[54][5] , \x[54][4] , \x[54][3] , \x[54][2] ,
         \x[54][1] , \x[54][0] , \x[53][15] , \x[53][14] , \x[53][13] ,
         \x[53][12] , \x[53][11] , \x[53][10] , \x[53][9] , \x[53][8] ,
         \x[53][7] , \x[53][6] , \x[53][5] , \x[53][4] , \x[53][3] ,
         \x[53][2] , \x[53][1] , \x[53][0] , \x[52][15] , \x[52][14] ,
         \x[52][13] , \x[52][12] , \x[52][11] , \x[52][10] , \x[52][9] ,
         \x[52][8] , \x[52][7] , \x[52][6] , \x[52][5] , \x[52][4] ,
         \x[52][3] , \x[52][2] , \x[52][1] , \x[52][0] , \x[51][15] ,
         \x[51][14] , \x[51][13] , \x[51][12] , \x[51][11] , \x[51][10] ,
         \x[51][9] , \x[51][8] , \x[51][7] , \x[51][6] , \x[51][5] ,
         \x[51][4] , \x[51][3] , \x[51][2] , \x[51][1] , \x[51][0] ,
         \x[50][15] , \x[50][14] , \x[50][13] , \x[50][12] , \x[50][11] ,
         \x[50][10] , \x[50][9] , \x[50][8] , \x[50][7] , \x[50][6] ,
         \x[50][5] , \x[50][4] , \x[50][3] , \x[50][2] , \x[50][1] ,
         \x[50][0] , \x[49][15] , \x[49][14] , \x[49][13] , \x[49][12] ,
         \x[49][11] , \x[49][10] , \x[49][9] , \x[49][8] , \x[49][7] ,
         \x[49][6] , \x[49][5] , \x[49][4] , \x[49][3] , \x[49][2] ,
         \x[49][1] , \x[49][0] , \x[48][15] , \x[48][14] , \x[48][13] ,
         \x[48][12] , \x[48][11] , \x[48][10] , \x[48][9] , \x[48][8] ,
         \x[48][7] , \x[48][6] , \x[48][5] , \x[48][4] , \x[48][3] ,
         \x[48][2] , \x[48][1] , \x[48][0] , \x[47][15] , \x[47][14] ,
         \x[47][13] , \x[47][12] , \x[47][11] , \x[47][10] , \x[47][9] ,
         \x[47][8] , \x[47][7] , \x[47][6] , \x[47][5] , \x[47][4] ,
         \x[47][3] , \x[47][2] , \x[47][1] , \x[47][0] , \x[46][15] ,
         \x[46][14] , \x[46][13] , \x[46][12] , \x[46][11] , \x[46][10] ,
         \x[46][9] , \x[46][8] , \x[46][7] , \x[46][6] , \x[46][5] ,
         \x[46][4] , \x[46][3] , \x[46][2] , \x[46][1] , \x[46][0] ,
         \x[45][15] , \x[45][14] , \x[45][13] , \x[45][12] , \x[45][11] ,
         \x[45][10] , \x[45][9] , \x[45][8] , \x[45][7] , \x[45][6] ,
         \x[45][5] , \x[45][4] , \x[45][3] , \x[45][2] , \x[45][1] ,
         \x[45][0] , \x[44][15] , \x[44][14] , \x[44][13] , \x[44][12] ,
         \x[44][11] , \x[44][10] , \x[44][9] , \x[44][8] , \x[44][7] ,
         \x[44][6] , \x[44][5] , \x[44][4] , \x[44][3] , \x[44][2] ,
         \x[44][1] , \x[44][0] , \x[43][15] , \x[43][14] , \x[43][13] ,
         \x[43][12] , \x[43][11] , \x[43][10] , \x[43][9] , \x[43][8] ,
         \x[43][7] , \x[43][6] , \x[43][5] , \x[43][4] , \x[43][3] ,
         \x[43][2] , \x[43][1] , \x[43][0] , \x[42][15] , \x[42][14] ,
         \x[42][13] , \x[42][12] , \x[42][11] , \x[42][10] , \x[42][9] ,
         \x[42][8] , \x[42][7] , \x[42][6] , \x[42][5] , \x[42][4] ,
         \x[42][3] , \x[42][2] , \x[42][1] , \x[42][0] , \x[41][15] ,
         \x[41][14] , \x[41][13] , \x[41][12] , \x[41][11] , \x[41][10] ,
         \x[41][9] , \x[41][8] , \x[41][7] , \x[41][6] , \x[41][5] ,
         \x[41][4] , \x[41][3] , \x[41][2] , \x[41][1] , \x[41][0] ,
         \x[40][15] , \x[40][14] , \x[40][13] , \x[40][12] , \x[40][11] ,
         \x[40][10] , \x[40][9] , \x[40][8] , \x[40][7] , \x[40][6] ,
         \x[40][5] , \x[40][4] , \x[40][3] , \x[40][2] , \x[40][1] ,
         \x[40][0] , \x[39][15] , \x[39][14] , \x[39][13] , \x[39][12] ,
         \x[39][11] , \x[39][10] , \x[39][9] , \x[39][8] , \x[39][7] ,
         \x[39][6] , \x[39][5] , \x[39][4] , \x[39][3] , \x[39][2] ,
         \x[39][1] , \x[39][0] , \x[38][15] , \x[38][14] , \x[38][13] ,
         \x[38][12] , \x[38][11] , \x[38][10] , \x[38][9] , \x[38][8] ,
         \x[38][7] , \x[38][6] , \x[38][5] , \x[38][4] , \x[38][3] ,
         \x[38][2] , \x[38][1] , \x[38][0] , \x[37][15] , \x[37][14] ,
         \x[37][13] , \x[37][12] , \x[37][11] , \x[37][10] , \x[37][9] ,
         \x[37][8] , \x[37][7] , \x[37][6] , \x[37][5] , \x[37][4] ,
         \x[37][3] , \x[37][2] , \x[37][1] , \x[37][0] , \x[36][15] ,
         \x[36][14] , \x[36][13] , \x[36][12] , \x[36][11] , \x[36][10] ,
         \x[36][9] , \x[36][8] , \x[36][7] , \x[36][6] , \x[36][5] ,
         \x[36][4] , \x[36][3] , \x[36][2] , \x[36][1] , \x[36][0] ,
         \x[35][15] , \x[35][14] , \x[35][13] , \x[35][12] , \x[35][11] ,
         \x[35][10] , \x[35][9] , \x[35][8] , \x[35][7] , \x[35][6] ,
         \x[35][5] , \x[35][4] , \x[35][3] , \x[35][2] , \x[35][1] ,
         \x[35][0] , \x[34][15] , \x[34][14] , \x[34][13] , \x[34][12] ,
         \x[34][11] , \x[34][10] , \x[34][9] , \x[34][8] , \x[34][7] ,
         \x[34][6] , \x[34][5] , \x[34][4] , \x[34][3] , \x[34][2] ,
         \x[34][1] , \x[34][0] , \x[33][15] , \x[33][14] , \x[33][13] ,
         \x[33][12] , \x[33][11] , \x[33][10] , \x[33][9] , \x[33][8] ,
         \x[33][7] , \x[33][6] , \x[33][5] , \x[33][4] , \x[33][3] ,
         \x[33][2] , \x[33][1] , \x[33][0] , \x[32][15] , \x[32][14] ,
         \x[32][13] , \x[32][12] , \x[32][11] , \x[32][10] , \x[32][9] ,
         \x[32][8] , \x[32][7] , \x[32][6] , \x[32][5] , \x[32][4] ,
         \x[32][3] , \x[32][2] , \x[32][1] , \x[32][0] , \x[31][15] ,
         \x[31][14] , \x[31][13] , \x[31][12] , \x[31][11] , \x[31][10] ,
         \x[31][9] , \x[31][8] , \x[31][7] , \x[31][6] , \x[31][5] ,
         \x[31][4] , \x[31][3] , \x[31][2] , \x[31][1] , \x[31][0] ,
         \x[30][15] , \x[30][14] , \x[30][13] , \x[30][12] , \x[30][11] ,
         \x[30][10] , \x[30][9] , \x[30][8] , \x[30][7] , \x[30][6] ,
         \x[30][5] , \x[30][4] , \x[30][3] , \x[30][2] , \x[30][1] ,
         \x[30][0] , \x[29][15] , \x[29][14] , \x[29][13] , \x[29][12] ,
         \x[29][11] , \x[29][10] , \x[29][9] , \x[29][8] , \x[29][7] ,
         \x[29][6] , \x[29][5] , \x[29][4] , \x[29][3] , \x[29][2] ,
         \x[29][1] , \x[29][0] , \x[28][15] , \x[28][14] , \x[28][13] ,
         \x[28][12] , \x[28][11] , \x[28][10] , \x[28][9] , \x[28][8] ,
         \x[28][7] , \x[28][6] , \x[28][5] , \x[28][4] , \x[28][3] ,
         \x[28][2] , \x[28][1] , \x[28][0] , \x[27][15] , \x[27][14] ,
         \x[27][13] , \x[27][12] , \x[27][11] , \x[27][10] , \x[27][9] ,
         \x[27][8] , \x[27][7] , \x[27][6] , \x[27][5] , \x[27][4] ,
         \x[27][3] , \x[27][2] , \x[27][1] , \x[27][0] , \x[26][15] ,
         \x[26][14] , \x[26][13] , \x[26][12] , \x[26][11] , \x[26][10] ,
         \x[26][9] , \x[26][8] , \x[26][7] , \x[26][6] , \x[26][5] ,
         \x[26][4] , \x[26][3] , \x[26][2] , \x[26][1] , \x[26][0] ,
         \x[25][15] , \x[25][14] , \x[25][13] , \x[25][12] , \x[25][11] ,
         \x[25][10] , \x[25][9] , \x[25][8] , \x[25][7] , \x[25][6] ,
         \x[25][5] , \x[25][4] , \x[25][3] , \x[25][2] , \x[25][1] ,
         \x[25][0] , \x[24][15] , \x[24][14] , \x[24][13] , \x[24][12] ,
         \x[24][11] , \x[24][10] , \x[24][9] , \x[24][8] , \x[24][7] ,
         \x[24][6] , \x[24][5] , \x[24][4] , \x[24][3] , \x[24][2] ,
         \x[24][1] , \x[24][0] , \x[23][15] , \x[23][14] , \x[23][13] ,
         \x[23][12] , \x[23][11] , \x[23][10] , \x[23][9] , \x[23][8] ,
         \x[23][7] , \x[23][6] , \x[23][5] , \x[23][4] , \x[23][3] ,
         \x[23][2] , \x[23][1] , \x[23][0] , \x[22][15] , \x[22][14] ,
         \x[22][13] , \x[22][12] , \x[22][11] , \x[22][10] , \x[22][9] ,
         \x[22][8] , \x[22][7] , \x[22][6] , \x[22][5] , \x[22][4] ,
         \x[22][3] , \x[22][2] , \x[22][1] , \x[22][0] , \x[21][15] ,
         \x[21][14] , \x[21][13] , \x[21][12] , \x[21][11] , \x[21][10] ,
         \x[21][9] , \x[21][8] , \x[21][7] , \x[21][6] , \x[21][5] ,
         \x[21][4] , \x[21][3] , \x[21][2] , \x[21][1] , \x[21][0] ,
         \x[20][15] , \x[20][14] , \x[20][13] , \x[20][12] , \x[20][11] ,
         \x[20][10] , \x[20][9] , \x[20][8] , \x[20][7] , \x[20][6] ,
         \x[20][5] , \x[20][4] , \x[20][3] , \x[20][2] , \x[20][1] ,
         \x[20][0] , \x[19][15] , \x[19][14] , \x[19][13] , \x[19][12] ,
         \x[19][11] , \x[19][10] , \x[19][9] , \x[19][8] , \x[19][7] ,
         \x[19][6] , \x[19][5] , \x[19][4] , \x[19][3] , \x[19][2] ,
         \x[19][1] , \x[19][0] , \x[18][15] , \x[18][14] , \x[18][13] ,
         \x[18][12] , \x[18][11] , \x[18][10] , \x[18][9] , \x[18][8] ,
         \x[18][7] , \x[18][6] , \x[18][5] , \x[18][4] , \x[18][3] ,
         \x[18][2] , \x[18][1] , \x[18][0] , \x[17][15] , \x[17][14] ,
         \x[17][13] , \x[17][12] , \x[17][11] , \x[17][10] , \x[17][9] ,
         \x[17][8] , \x[17][7] , \x[17][6] , \x[17][5] , \x[17][4] ,
         \x[17][3] , \x[17][2] , \x[17][1] , \x[17][0] , \x[16][15] ,
         \x[16][14] , \x[16][13] , \x[16][12] , \x[16][11] , \x[16][10] ,
         \x[16][9] , \x[16][8] , \x[16][7] , \x[16][6] , \x[16][5] ,
         \x[16][4] , \x[16][3] , \x[16][2] , \x[16][1] , \x[16][0] ,
         \x[15][15] , \x[15][14] , \x[15][13] , \x[15][12] , \x[15][11] ,
         \x[15][10] , \x[15][9] , \x[15][8] , \x[15][7] , \x[15][6] ,
         \x[15][5] , \x[15][4] , \x[15][3] , \x[15][2] , \x[15][1] ,
         \x[15][0] , \x[14][15] , \x[14][14] , \x[14][13] , \x[14][12] ,
         \x[14][11] , \x[14][10] , \x[14][9] , \x[14][8] , \x[14][7] ,
         \x[14][6] , \x[14][5] , \x[14][4] , \x[14][3] , \x[14][2] ,
         \x[14][1] , \x[14][0] , \x[13][15] , \x[13][14] , \x[13][13] ,
         \x[13][12] , \x[13][11] , \x[13][10] , \x[13][9] , \x[13][8] ,
         \x[13][7] , \x[13][6] , \x[13][5] , \x[13][4] , \x[13][3] ,
         \x[13][2] , \x[13][1] , \x[13][0] , \x[12][15] , \x[12][14] ,
         \x[12][13] , \x[12][12] , \x[12][11] , \x[12][10] , \x[12][9] ,
         \x[12][8] , \x[12][7] , \x[12][6] , \x[12][5] , \x[12][4] ,
         \x[12][3] , \x[12][2] , \x[12][1] , \x[12][0] , \x[11][15] ,
         \x[11][14] , \x[11][13] , \x[11][12] , \x[11][11] , \x[11][10] ,
         \x[11][9] , \x[11][8] , \x[11][7] , \x[11][6] , \x[11][5] ,
         \x[11][4] , \x[11][3] , \x[11][2] , \x[11][1] , \x[11][0] ,
         \x[10][15] , \x[10][14] , \x[10][13] , \x[10][12] , \x[10][11] ,
         \x[10][10] , \x[10][9] , \x[10][8] , \x[10][7] , \x[10][6] ,
         \x[10][5] , \x[10][4] , \x[10][3] , \x[10][2] , \x[10][1] ,
         \x[10][0] , \x[9][15] , \x[9][14] , \x[9][13] , \x[9][12] ,
         \x[9][11] , \x[9][10] , \x[9][9] , \x[9][8] , \x[9][7] , \x[9][6] ,
         \x[9][5] , \x[9][4] , \x[9][3] , \x[9][2] , \x[9][1] , \x[9][0] ,
         \x[8][15] , \x[8][14] , \x[8][13] , \x[8][12] , \x[8][11] ,
         \x[8][10] , \x[8][9] , \x[8][8] , \x[8][7] , \x[8][6] , \x[8][5] ,
         \x[8][4] , \x[8][3] , \x[8][2] , \x[8][1] , \x[8][0] , \x[7][15] ,
         \x[7][14] , \x[7][13] , \x[7][12] , \x[7][11] , \x[7][10] , \x[7][9] ,
         \x[7][8] , \x[7][7] , \x[7][6] , \x[7][5] , \x[7][4] , \x[7][3] ,
         \x[7][2] , \x[7][1] , \x[7][0] , \x[6][15] , \x[6][14] , \x[6][13] ,
         \x[6][12] , \x[6][11] , \x[6][10] , \x[6][9] , \x[6][8] , \x[6][7] ,
         \x[6][6] , \x[6][5] , \x[6][4] , \x[6][3] , \x[6][2] , \x[6][1] ,
         \x[6][0] , \x[5][15] , \x[5][14] , \x[5][13] , \x[5][12] , \x[5][11] ,
         \x[5][10] , \x[5][9] , \x[5][8] , \x[5][7] , \x[5][6] , \x[5][5] ,
         \x[5][4] , \x[5][3] , \x[5][2] , \x[5][1] , \x[5][0] , \x[4][15] ,
         \x[4][14] , \x[4][13] , \x[4][12] , \x[4][11] , \x[4][10] , \x[4][9] ,
         \x[4][8] , \x[4][7] , \x[4][6] , \x[4][5] , \x[4][4] , \x[4][3] ,
         \x[4][2] , \x[4][1] , \x[4][0] , \x[3][15] , \x[3][14] , \x[3][13] ,
         \x[3][12] , \x[3][11] , \x[3][10] , \x[3][9] , \x[3][8] , \x[3][7] ,
         \x[3][6] , \x[3][5] , \x[3][4] , \x[3][3] , \x[3][2] , \x[3][1] ,
         \x[3][0] , \x[2][15] , \x[2][14] , \x[2][13] , \x[2][12] , \x[2][11] ,
         \x[2][10] , \x[2][9] , \x[2][8] , \x[2][7] , \x[2][6] , \x[2][5] ,
         \x[2][4] , \x[2][3] , \x[2][2] , \x[2][1] , \x[2][0] , \x[1][15] ,
         \x[1][14] , \x[1][13] , \x[1][12] , \x[1][11] , \x[1][10] , \x[1][9] ,
         \x[1][8] , \x[1][7] , \x[1][6] , \x[1][5] , \x[1][4] , \x[1][3] ,
         \x[1][2] , \x[1][1] , \x[1][0] , \x[0][15] , \x[0][14] , \x[0][13] ,
         \x[0][12] , \x[0][11] , \x[0][10] , \x[0][9] , \x[0][8] , \x[0][7] ,
         \x[0][6] , \x[0][5] , \x[0][4] , \x[0][3] , \x[0][2] , \x[0][1] ,
         \x[0][0] , \LUT[24][15] , \LUT[24][14] , \LUT[24][13] , \LUT[24][12] ,
         \LUT[24][11] , \LUT[24][10] , \LUT[24][9] , \LUT[24][8] ,
         \LUT[24][7] , \LUT[24][6] , \LUT[24][5] , \LUT[24][4] , \LUT[24][3] ,
         \LUT[24][2] , \LUT[24][1] , \LUT[24][0] , \LUT[23][15] ,
         \LUT[23][14] , \LUT[23][13] , \LUT[23][12] , \LUT[23][11] ,
         \LUT[23][10] , \LUT[23][9] , \LUT[23][8] , \LUT[23][7] , \LUT[23][6] ,
         \LUT[23][5] , \LUT[23][4] , \LUT[23][3] , \LUT[23][2] , \LUT[23][1] ,
         \LUT[23][0] , \LUT[22][15] , \LUT[22][14] , \LUT[22][13] ,
         \LUT[22][12] , \LUT[22][11] , \LUT[22][10] , \LUT[22][9] ,
         \LUT[22][8] , \LUT[22][7] , \LUT[22][6] , \LUT[22][5] , \LUT[22][4] ,
         \LUT[22][3] , \LUT[22][2] , \LUT[22][1] , \LUT[22][0] , \LUT[21][15] ,
         \LUT[21][14] , \LUT[21][13] , \LUT[21][12] , \LUT[21][11] ,
         \LUT[21][10] , \LUT[21][9] , \LUT[21][8] , \LUT[21][7] , \LUT[21][6] ,
         \LUT[21][5] , \LUT[21][4] , \LUT[21][3] , \LUT[21][2] , \LUT[21][1] ,
         \LUT[21][0] , \LUT[20][15] , \LUT[20][14] , \LUT[20][13] ,
         \LUT[20][12] , \LUT[20][11] , \LUT[20][10] , \LUT[20][9] ,
         \LUT[20][8] , \LUT[20][7] , \LUT[20][6] , \LUT[20][5] , \LUT[20][4] ,
         \LUT[20][3] , \LUT[20][2] , \LUT[20][1] , \LUT[20][0] , \LUT[19][15] ,
         \LUT[19][14] , \LUT[19][13] , \LUT[19][12] , \LUT[19][11] ,
         \LUT[19][10] , \LUT[19][9] , \LUT[19][8] , \LUT[19][7] , \LUT[19][6] ,
         \LUT[19][5] , \LUT[19][4] , \LUT[19][3] , \LUT[19][2] , \LUT[19][1] ,
         \LUT[19][0] , \LUT[18][15] , \LUT[18][14] , \LUT[18][13] ,
         \LUT[18][12] , \LUT[18][11] , \LUT[18][10] , \LUT[18][9] ,
         \LUT[18][8] , \LUT[18][7] , \LUT[18][6] , \LUT[18][5] , \LUT[18][4] ,
         \LUT[18][3] , \LUT[18][2] , \LUT[18][1] , \LUT[18][0] , \LUT[17][15] ,
         \LUT[17][14] , \LUT[17][13] , \LUT[17][12] , \LUT[17][11] ,
         \LUT[17][10] , \LUT[17][9] , \LUT[17][8] , \LUT[17][7] , \LUT[17][6] ,
         \LUT[17][5] , \LUT[17][4] , \LUT[17][3] , \LUT[17][2] , \LUT[17][1] ,
         \LUT[17][0] , \LUT[16][15] , \LUT[16][14] , \LUT[16][13] ,
         \LUT[16][12] , \LUT[16][11] , \LUT[16][10] , \LUT[16][9] ,
         \LUT[16][8] , \LUT[16][7] , \LUT[16][6] , \LUT[16][5] , \LUT[16][4] ,
         \LUT[16][3] , \LUT[16][2] , \LUT[16][1] , \LUT[16][0] , \LUT[15][15] ,
         \LUT[15][14] , \LUT[15][13] , \LUT[15][12] , \LUT[15][11] ,
         \LUT[15][10] , \LUT[15][9] , \LUT[15][8] , \LUT[15][7] , \LUT[15][6] ,
         \LUT[15][5] , \LUT[15][4] , \LUT[15][3] , \LUT[15][2] , \LUT[15][1] ,
         \LUT[15][0] , \LUT[14][15] , \LUT[14][14] , \LUT[14][13] ,
         \LUT[14][12] , \LUT[14][11] , \LUT[14][10] , \LUT[14][9] ,
         \LUT[14][8] , \LUT[14][7] , \LUT[14][6] , \LUT[14][5] , \LUT[14][4] ,
         \LUT[14][3] , \LUT[14][2] , \LUT[14][1] , \LUT[14][0] , \LUT[13][15] ,
         \LUT[13][14] , \LUT[13][13] , \LUT[13][12] , \LUT[13][11] ,
         \LUT[13][10] , \LUT[13][9] , \LUT[13][8] , \LUT[13][7] , \LUT[13][6] ,
         \LUT[13][5] , \LUT[13][4] , \LUT[13][3] , \LUT[13][2] , \LUT[13][1] ,
         \LUT[13][0] , \LUT[12][15] , \LUT[12][14] , \LUT[12][13] ,
         \LUT[12][12] , \LUT[12][11] , \LUT[12][10] , \LUT[12][9] ,
         \LUT[12][8] , \LUT[12][7] , \LUT[12][6] , \LUT[12][5] , \LUT[12][4] ,
         \LUT[12][3] , \LUT[12][2] , \LUT[12][1] , \LUT[12][0] , \LUT[11][15] ,
         \LUT[11][14] , \LUT[11][13] , \LUT[11][12] , \LUT[11][11] ,
         \LUT[11][10] , \LUT[11][9] , \LUT[11][8] , \LUT[11][7] , \LUT[11][6] ,
         \LUT[11][5] , \LUT[11][4] , \LUT[11][3] , \LUT[11][2] , \LUT[11][1] ,
         \LUT[11][0] , \LUT[10][15] , \LUT[10][14] , \LUT[10][13] ,
         \LUT[10][12] , \LUT[10][11] , \LUT[10][10] , \LUT[10][9] ,
         \LUT[10][8] , \LUT[10][7] , \LUT[10][6] , \LUT[10][5] , \LUT[10][4] ,
         \LUT[10][3] , \LUT[10][2] , \LUT[10][1] , \LUT[10][0] , \LUT[9][15] ,
         \LUT[9][14] , \LUT[9][13] , \LUT[9][12] , \LUT[9][11] , \LUT[9][10] ,
         \LUT[9][9] , \LUT[9][8] , \LUT[9][7] , \LUT[9][6] , \LUT[9][5] ,
         \LUT[9][4] , \LUT[9][3] , \LUT[9][2] , \LUT[9][1] , \LUT[9][0] ,
         \LUT[8][15] , \LUT[8][14] , \LUT[8][13] , \LUT[8][12] , \LUT[8][11] ,
         \LUT[8][10] , \LUT[8][9] , \LUT[8][8] , \LUT[8][7] , \LUT[8][6] ,
         \LUT[8][5] , \LUT[8][4] , \LUT[8][3] , \LUT[8][2] , \LUT[8][1] ,
         \LUT[8][0] , \LUT[7][15] , \LUT[7][14] , \LUT[7][13] , \LUT[7][12] ,
         \LUT[7][11] , \LUT[7][10] , \LUT[7][9] , \LUT[7][8] , \LUT[7][7] ,
         \LUT[7][6] , \LUT[7][5] , \LUT[7][4] , \LUT[7][3] , \LUT[7][2] ,
         \LUT[7][1] , \LUT[7][0] , \LUT[6][15] , \LUT[6][14] , \LUT[6][13] ,
         \LUT[6][12] , \LUT[6][11] , \LUT[6][10] , \LUT[6][9] , \LUT[6][8] ,
         \LUT[6][7] , \LUT[6][6] , \LUT[6][5] , \LUT[6][4] , \LUT[6][3] ,
         \LUT[6][2] , \LUT[6][1] , \LUT[6][0] , \LUT[5][15] , \LUT[5][14] ,
         \LUT[5][13] , \LUT[5][12] , \LUT[5][11] , \LUT[5][10] , \LUT[5][9] ,
         \LUT[5][8] , \LUT[5][7] , \LUT[5][6] , \LUT[5][5] , \LUT[5][4] ,
         \LUT[5][3] , \LUT[5][2] , \LUT[5][1] , \LUT[5][0] , \LUT[4][15] ,
         \LUT[4][14] , \LUT[4][13] , \LUT[4][12] , \LUT[4][11] , \LUT[4][10] ,
         \LUT[4][9] , \LUT[4][8] , \LUT[4][7] , \LUT[4][6] , \LUT[4][5] ,
         \LUT[4][4] , \LUT[4][3] , \LUT[4][2] , \LUT[4][1] , \LUT[4][0] ,
         \LUT[3][15] , \LUT[3][14] , \LUT[3][13] , \LUT[3][12] , \LUT[3][11] ,
         \LUT[3][10] , \LUT[3][9] , \LUT[3][8] , \LUT[3][7] , \LUT[3][6] ,
         \LUT[3][5] , \LUT[3][4] , \LUT[3][3] , \LUT[3][2] , \LUT[3][1] ,
         \LUT[3][0] , \LUT[2][15] , \LUT[2][14] , \LUT[2][13] , \LUT[2][12] ,
         \LUT[2][11] , \LUT[2][10] , \LUT[2][9] , \LUT[2][8] , \LUT[2][7] ,
         \LUT[2][6] , \LUT[2][5] , \LUT[2][4] , \LUT[2][3] , \LUT[2][2] ,
         \LUT[2][1] , \LUT[2][0] , \LUT[1][15] , \LUT[1][14] , \LUT[1][13] ,
         \LUT[1][12] , \LUT[1][11] , \LUT[1][10] , \LUT[1][9] , \LUT[1][8] ,
         \LUT[1][7] , \LUT[1][6] , \LUT[1][5] , \LUT[1][4] , \LUT[1][3] ,
         \LUT[1][2] , \LUT[1][1] , \LUT[1][0] , \LUT[0][15] , \LUT[0][14] ,
         \LUT[0][13] , \LUT[0][12] , \LUT[0][11] , \LUT[0][10] , \LUT[0][9] ,
         \LUT[0][8] , \LUT[0][7] , \LUT[0][6] , \LUT[0][5] , \LUT[0][4] ,
         \LUT[0][3] , \LUT[0][2] , \LUT[0][1] , \LUT[0][0] , \LUT[56][15] ,
         \LUT[56][14] , \LUT[56][13] , \LUT[56][12] , \LUT[56][11] ,
         \LUT[56][10] , \LUT[56][9] , \LUT[56][8] , \LUT[56][7] , \LUT[56][6] ,
         \LUT[56][5] , \LUT[56][4] , \LUT[56][3] , \LUT[56][2] , \LUT[56][1] ,
         \LUT[56][0] , \LUT[55][15] , \LUT[55][14] , \LUT[55][13] ,
         \LUT[55][12] , \LUT[55][11] , \LUT[55][10] , \LUT[55][9] ,
         \LUT[55][8] , \LUT[55][7] , \LUT[55][6] , \LUT[55][5] , \LUT[55][4] ,
         \LUT[55][3] , \LUT[55][2] , \LUT[55][1] , \LUT[55][0] , \LUT[54][15] ,
         \LUT[54][14] , \LUT[54][13] , \LUT[54][12] , \LUT[54][11] ,
         \LUT[54][10] , \LUT[54][9] , \LUT[54][8] , \LUT[54][7] , \LUT[54][6] ,
         \LUT[54][5] , \LUT[54][4] , \LUT[54][3] , \LUT[54][2] , \LUT[54][1] ,
         \LUT[54][0] , \LUT[53][15] , \LUT[53][14] , \LUT[53][13] ,
         \LUT[53][12] , \LUT[53][11] , \LUT[53][10] , \LUT[53][9] ,
         \LUT[53][8] , \LUT[53][7] , \LUT[53][6] , \LUT[53][5] , \LUT[53][4] ,
         \LUT[53][3] , \LUT[53][2] , \LUT[53][1] , \LUT[53][0] , \LUT[52][15] ,
         \LUT[52][14] , \LUT[52][13] , \LUT[52][12] , \LUT[52][11] ,
         \LUT[52][10] , \LUT[52][9] , \LUT[52][8] , \LUT[52][7] , \LUT[52][6] ,
         \LUT[52][5] , \LUT[52][4] , \LUT[52][3] , \LUT[52][2] , \LUT[52][1] ,
         \LUT[52][0] , \LUT[51][15] , \LUT[51][14] , \LUT[51][13] ,
         \LUT[51][12] , \LUT[51][11] , \LUT[51][10] , \LUT[51][9] ,
         \LUT[51][8] , \LUT[51][7] , \LUT[51][6] , \LUT[51][5] , \LUT[51][4] ,
         \LUT[51][3] , \LUT[51][2] , \LUT[51][1] , \LUT[51][0] , \LUT[50][15] ,
         \LUT[50][14] , \LUT[50][13] , \LUT[50][12] , \LUT[50][11] ,
         \LUT[50][10] , \LUT[50][9] , \LUT[50][8] , \LUT[50][7] , \LUT[50][6] ,
         \LUT[50][5] , \LUT[50][4] , \LUT[50][3] , \LUT[50][2] , \LUT[50][1] ,
         \LUT[50][0] , \LUT[49][15] , \LUT[49][14] , \LUT[49][13] ,
         \LUT[49][12] , \LUT[49][11] , \LUT[49][10] , \LUT[49][9] ,
         \LUT[49][8] , \LUT[49][7] , \LUT[49][6] , \LUT[49][5] , \LUT[49][4] ,
         \LUT[49][3] , \LUT[49][2] , \LUT[49][1] , \LUT[49][0] , \LUT[48][15] ,
         \LUT[48][14] , \LUT[48][13] , \LUT[48][12] , \LUT[48][11] ,
         \LUT[48][10] , \LUT[48][9] , \LUT[48][8] , \LUT[48][7] , \LUT[48][6] ,
         \LUT[48][5] , \LUT[48][4] , \LUT[48][3] , \LUT[48][2] , \LUT[48][1] ,
         \LUT[48][0] , \LUT[47][15] , \LUT[47][14] , \LUT[47][13] ,
         \LUT[47][12] , \LUT[47][11] , \LUT[47][10] , \LUT[47][9] ,
         \LUT[47][8] , \LUT[47][7] , \LUT[47][6] , \LUT[47][5] , \LUT[47][4] ,
         \LUT[47][3] , \LUT[47][2] , \LUT[47][1] , \LUT[47][0] , \LUT[46][15] ,
         \LUT[46][14] , \LUT[46][13] , \LUT[46][12] , \LUT[46][11] ,
         \LUT[46][10] , \LUT[46][9] , \LUT[46][8] , \LUT[46][7] , \LUT[46][6] ,
         \LUT[46][5] , \LUT[46][4] , \LUT[46][3] , \LUT[46][2] , \LUT[46][1] ,
         \LUT[46][0] , \LUT[45][15] , \LUT[45][14] , \LUT[45][13] ,
         \LUT[45][12] , \LUT[45][11] , \LUT[45][10] , \LUT[45][9] ,
         \LUT[45][8] , \LUT[45][7] , \LUT[45][6] , \LUT[45][5] , \LUT[45][4] ,
         \LUT[45][3] , \LUT[45][2] , \LUT[45][1] , \LUT[45][0] , \LUT[44][15] ,
         \LUT[44][14] , \LUT[44][13] , \LUT[44][12] , \LUT[44][11] ,
         \LUT[44][10] , \LUT[44][9] , \LUT[44][8] , \LUT[44][7] , \LUT[44][6] ,
         \LUT[44][5] , \LUT[44][4] , \LUT[44][3] , \LUT[44][2] , \LUT[44][1] ,
         \LUT[44][0] , \LUT[43][15] , \LUT[43][14] , \LUT[43][13] ,
         \LUT[43][12] , \LUT[43][11] , \LUT[43][10] , \LUT[43][9] ,
         \LUT[43][8] , \LUT[43][7] , \LUT[43][6] , \LUT[43][5] , \LUT[43][4] ,
         \LUT[43][3] , \LUT[43][2] , \LUT[43][1] , \LUT[43][0] , \LUT[42][15] ,
         \LUT[42][14] , \LUT[42][13] , \LUT[42][12] , \LUT[42][11] ,
         \LUT[42][10] , \LUT[42][9] , \LUT[42][8] , \LUT[42][7] , \LUT[42][6] ,
         \LUT[42][5] , \LUT[42][4] , \LUT[42][3] , \LUT[42][2] , \LUT[42][1] ,
         \LUT[42][0] , \LUT[41][15] , \LUT[41][14] , \LUT[41][13] ,
         \LUT[41][12] , \LUT[41][11] , \LUT[41][10] , \LUT[41][9] ,
         \LUT[41][8] , \LUT[41][7] , \LUT[41][6] , \LUT[41][5] , \LUT[41][4] ,
         \LUT[41][3] , \LUT[41][2] , \LUT[41][1] , \LUT[41][0] , \LUT[40][15] ,
         \LUT[40][14] , \LUT[40][13] , \LUT[40][12] , \LUT[40][11] ,
         \LUT[40][10] , \LUT[40][9] , \LUT[40][8] , \LUT[40][7] , \LUT[40][6] ,
         \LUT[40][5] , \LUT[40][4] , \LUT[40][3] , \LUT[40][2] , \LUT[40][1] ,
         \LUT[40][0] , \LUT[39][15] , \LUT[39][14] , \LUT[39][13] ,
         \LUT[39][12] , \LUT[39][11] , \LUT[39][10] , \LUT[39][9] ,
         \LUT[39][8] , \LUT[39][7] , \LUT[39][6] , \LUT[39][5] , \LUT[39][4] ,
         \LUT[39][3] , \LUT[39][2] , \LUT[39][1] , \LUT[39][0] , \LUT[38][15] ,
         \LUT[38][14] , \LUT[38][13] , \LUT[38][12] , \LUT[38][11] ,
         \LUT[38][10] , \LUT[38][9] , \LUT[38][8] , \LUT[38][7] , \LUT[38][6] ,
         \LUT[38][5] , \LUT[38][4] , \LUT[38][3] , \LUT[38][2] , \LUT[38][1] ,
         \LUT[38][0] , \LUT[37][15] , \LUT[37][14] , \LUT[37][13] ,
         \LUT[37][12] , \LUT[37][11] , \LUT[37][10] , \LUT[37][9] ,
         \LUT[37][8] , \LUT[37][7] , \LUT[37][6] , \LUT[37][5] , \LUT[37][4] ,
         \LUT[37][3] , \LUT[37][2] , \LUT[37][1] , \LUT[37][0] , \LUT[36][15] ,
         \LUT[36][14] , \LUT[36][13] , \LUT[36][12] , \LUT[36][11] ,
         \LUT[36][10] , \LUT[36][9] , \LUT[36][8] , \LUT[36][7] , \LUT[36][6] ,
         \LUT[36][5] , \LUT[36][4] , \LUT[36][3] , \LUT[36][2] , \LUT[36][1] ,
         \LUT[36][0] , \LUT[35][15] , \LUT[35][14] , \LUT[35][13] ,
         \LUT[35][12] , \LUT[35][11] , \LUT[35][10] , \LUT[35][9] ,
         \LUT[35][8] , \LUT[35][7] , \LUT[35][6] , \LUT[35][5] , \LUT[35][4] ,
         \LUT[35][3] , \LUT[35][2] , \LUT[35][1] , \LUT[35][0] , \LUT[34][15] ,
         \LUT[34][14] , \LUT[34][13] , \LUT[34][12] , \LUT[34][11] ,
         \LUT[34][10] , \LUT[34][9] , \LUT[34][8] , \LUT[34][7] , \LUT[34][6] ,
         \LUT[34][5] , \LUT[34][4] , \LUT[34][3] , \LUT[34][2] , \LUT[34][1] ,
         \LUT[34][0] , \LUT[33][15] , \LUT[33][14] , \LUT[33][13] ,
         \LUT[33][12] , \LUT[33][11] , \LUT[33][10] , \LUT[33][9] ,
         \LUT[33][8] , \LUT[33][7] , \LUT[33][6] , \LUT[33][5] , \LUT[33][4] ,
         \LUT[33][3] , \LUT[33][2] , \LUT[33][1] , \LUT[33][0] , \LUT[32][15] ,
         \LUT[32][14] , \LUT[32][13] , \LUT[32][12] , \LUT[32][11] ,
         \LUT[32][10] , \LUT[32][9] , \LUT[32][8] , \LUT[32][7] , \LUT[32][6] ,
         \LUT[32][5] , \LUT[32][4] , \LUT[32][3] , \LUT[32][2] , \LUT[32][1] ,
         \LUT[32][0] , \LUT[31][15] , \LUT[31][14] , \LUT[31][13] ,
         \LUT[31][12] , \LUT[31][11] , \LUT[31][10] , \LUT[31][9] ,
         \LUT[31][8] , \LUT[31][7] , \LUT[31][6] , \LUT[31][5] , \LUT[31][4] ,
         \LUT[31][3] , \LUT[31][2] , \LUT[31][1] , \LUT[31][0] , \LUT[30][15] ,
         \LUT[30][14] , \LUT[30][13] , \LUT[30][12] , \LUT[30][11] ,
         \LUT[30][10] , \LUT[30][9] , \LUT[30][8] , \LUT[30][7] , \LUT[30][6] ,
         \LUT[30][5] , \LUT[30][4] , \LUT[30][3] , \LUT[30][2] , \LUT[30][1] ,
         \LUT[30][0] , \LUT[29][15] , \LUT[29][14] , \LUT[29][13] ,
         \LUT[29][12] , \LUT[29][11] , \LUT[29][10] , \LUT[29][9] ,
         \LUT[29][8] , \LUT[29][7] , \LUT[29][6] , \LUT[29][5] , \LUT[29][4] ,
         \LUT[29][3] , \LUT[29][2] , \LUT[29][1] , \LUT[29][0] , \LUT[28][15] ,
         \LUT[28][14] , \LUT[28][13] , \LUT[28][12] , \LUT[28][11] ,
         \LUT[28][10] , \LUT[28][9] , \LUT[28][8] , \LUT[28][7] , \LUT[28][6] ,
         \LUT[28][5] , \LUT[28][4] , \LUT[28][3] , \LUT[28][2] , \LUT[28][1] ,
         \LUT[28][0] , \LUT[27][15] , \LUT[27][14] , \LUT[27][13] ,
         \LUT[27][12] , \LUT[27][11] , \LUT[27][10] , \LUT[27][9] ,
         \LUT[27][8] , \LUT[27][7] , \LUT[27][6] , \LUT[27][5] , \LUT[27][4] ,
         \LUT[27][3] , \LUT[27][2] , \LUT[27][1] , \LUT[27][0] , \LUT[26][15] ,
         \LUT[26][14] , \LUT[26][13] , \LUT[26][12] , \LUT[26][11] ,
         \LUT[26][10] , \LUT[26][9] , \LUT[26][8] , \LUT[26][7] , \LUT[26][6] ,
         \LUT[26][5] , \LUT[26][4] , \LUT[26][3] , \LUT[26][2] , \LUT[26][1] ,
         \LUT[26][0] , \LUT[25][15] , \LUT[25][14] , \LUT[25][13] ,
         \LUT[25][12] , \LUT[25][11] , \LUT[25][10] , \LUT[25][9] ,
         \LUT[25][8] , \LUT[25][7] , \LUT[25][6] , \LUT[25][5] , \LUT[25][4] ,
         \LUT[25][3] , \LUT[25][2] , \LUT[25][1] , \LUT[25][0] , \LUT[88][15] ,
         \LUT[88][14] , \LUT[88][13] , \LUT[88][12] , \LUT[88][11] ,
         \LUT[88][10] , \LUT[88][9] , \LUT[88][8] , \LUT[88][7] , \LUT[88][6] ,
         \LUT[88][5] , \LUT[88][4] , \LUT[88][3] , \LUT[88][2] , \LUT[88][1] ,
         \LUT[88][0] , \LUT[87][15] , \LUT[87][14] , \LUT[87][13] ,
         \LUT[87][12] , \LUT[87][11] , \LUT[87][10] , \LUT[87][9] ,
         \LUT[87][8] , \LUT[87][7] , \LUT[87][6] , \LUT[87][5] , \LUT[87][4] ,
         \LUT[87][3] , \LUT[87][2] , \LUT[87][1] , \LUT[87][0] , \LUT[86][15] ,
         \LUT[86][14] , \LUT[86][13] , \LUT[86][12] , \LUT[86][11] ,
         \LUT[86][10] , \LUT[86][9] , \LUT[86][8] , \LUT[86][7] , \LUT[86][6] ,
         \LUT[86][5] , \LUT[86][4] , \LUT[86][3] , \LUT[86][2] , \LUT[86][1] ,
         \LUT[86][0] , \LUT[85][15] , \LUT[85][14] , \LUT[85][13] ,
         \LUT[85][12] , \LUT[85][11] , \LUT[85][10] , \LUT[85][9] ,
         \LUT[85][8] , \LUT[85][7] , \LUT[85][6] , \LUT[85][5] , \LUT[85][4] ,
         \LUT[85][3] , \LUT[85][2] , \LUT[85][1] , \LUT[85][0] , \LUT[84][15] ,
         \LUT[84][14] , \LUT[84][13] , \LUT[84][12] , \LUT[84][11] ,
         \LUT[84][10] , \LUT[84][9] , \LUT[84][8] , \LUT[84][7] , \LUT[84][6] ,
         \LUT[84][5] , \LUT[84][4] , \LUT[84][3] , \LUT[84][2] , \LUT[84][1] ,
         \LUT[84][0] , \LUT[83][15] , \LUT[83][14] , \LUT[83][13] ,
         \LUT[83][12] , \LUT[83][11] , \LUT[83][10] , \LUT[83][9] ,
         \LUT[83][8] , \LUT[83][7] , \LUT[83][6] , \LUT[83][5] , \LUT[83][4] ,
         \LUT[83][3] , \LUT[83][2] , \LUT[83][1] , \LUT[83][0] , \LUT[82][15] ,
         \LUT[82][14] , \LUT[82][13] , \LUT[82][12] , \LUT[82][11] ,
         \LUT[82][10] , \LUT[82][9] , \LUT[82][8] , \LUT[82][7] , \LUT[82][6] ,
         \LUT[82][5] , \LUT[82][4] , \LUT[82][3] , \LUT[82][2] , \LUT[82][1] ,
         \LUT[82][0] , \LUT[81][15] , \LUT[81][14] , \LUT[81][13] ,
         \LUT[81][12] , \LUT[81][11] , \LUT[81][10] , \LUT[81][9] ,
         \LUT[81][8] , \LUT[81][7] , \LUT[81][6] , \LUT[81][5] , \LUT[81][4] ,
         \LUT[81][3] , \LUT[81][2] , \LUT[81][1] , \LUT[81][0] , \LUT[80][15] ,
         \LUT[80][14] , \LUT[80][13] , \LUT[80][12] , \LUT[80][11] ,
         \LUT[80][10] , \LUT[80][9] , \LUT[80][8] , \LUT[80][7] , \LUT[80][6] ,
         \LUT[80][5] , \LUT[80][4] , \LUT[80][3] , \LUT[80][2] , \LUT[80][1] ,
         \LUT[80][0] , \LUT[79][15] , \LUT[79][14] , \LUT[79][13] ,
         \LUT[79][12] , \LUT[79][11] , \LUT[79][10] , \LUT[79][9] ,
         \LUT[79][8] , \LUT[79][7] , \LUT[79][6] , \LUT[79][5] , \LUT[79][4] ,
         \LUT[79][3] , \LUT[79][2] , \LUT[79][1] , \LUT[79][0] , \LUT[78][15] ,
         \LUT[78][14] , \LUT[78][13] , \LUT[78][12] , \LUT[78][11] ,
         \LUT[78][10] , \LUT[78][9] , \LUT[78][8] , \LUT[78][7] , \LUT[78][6] ,
         \LUT[78][5] , \LUT[78][4] , \LUT[78][3] , \LUT[78][2] , \LUT[78][1] ,
         \LUT[78][0] , \LUT[77][15] , \LUT[77][14] , \LUT[77][13] ,
         \LUT[77][12] , \LUT[77][11] , \LUT[77][10] , \LUT[77][9] ,
         \LUT[77][8] , \LUT[77][7] , \LUT[77][6] , \LUT[77][5] , \LUT[77][4] ,
         \LUT[77][3] , \LUT[77][2] , \LUT[77][1] , \LUT[77][0] , \LUT[76][15] ,
         \LUT[76][14] , \LUT[76][13] , \LUT[76][12] , \LUT[76][11] ,
         \LUT[76][10] , \LUT[76][9] , \LUT[76][8] , \LUT[76][7] , \LUT[76][6] ,
         \LUT[76][5] , \LUT[76][4] , \LUT[76][3] , \LUT[76][2] , \LUT[76][1] ,
         \LUT[76][0] , \LUT[75][15] , \LUT[75][14] , \LUT[75][13] ,
         \LUT[75][12] , \LUT[75][11] , \LUT[75][10] , \LUT[75][9] ,
         \LUT[75][8] , \LUT[75][7] , \LUT[75][6] , \LUT[75][5] , \LUT[75][4] ,
         \LUT[75][3] , \LUT[75][2] , \LUT[75][1] , \LUT[75][0] , \LUT[74][15] ,
         \LUT[74][14] , \LUT[74][13] , \LUT[74][12] , \LUT[74][11] ,
         \LUT[74][10] , \LUT[74][9] , \LUT[74][8] , \LUT[74][7] , \LUT[74][6] ,
         \LUT[74][5] , \LUT[74][4] , \LUT[74][3] , \LUT[74][2] , \LUT[74][1] ,
         \LUT[74][0] , \LUT[73][15] , \LUT[73][14] , \LUT[73][13] ,
         \LUT[73][12] , \LUT[73][11] , \LUT[73][10] , \LUT[73][9] ,
         \LUT[73][8] , \LUT[73][7] , \LUT[73][6] , \LUT[73][5] , \LUT[73][4] ,
         \LUT[73][3] , \LUT[73][2] , \LUT[73][1] , \LUT[73][0] , \LUT[72][15] ,
         \LUT[72][14] , \LUT[72][13] , \LUT[72][12] , \LUT[72][11] ,
         \LUT[72][10] , \LUT[72][9] , \LUT[72][8] , \LUT[72][7] , \LUT[72][6] ,
         \LUT[72][5] , \LUT[72][4] , \LUT[72][3] , \LUT[72][2] , \LUT[72][1] ,
         \LUT[72][0] , \LUT[71][15] , \LUT[71][14] , \LUT[71][13] ,
         \LUT[71][12] , \LUT[71][11] , \LUT[71][10] , \LUT[71][9] ,
         \LUT[71][8] , \LUT[71][7] , \LUT[71][6] , \LUT[71][5] , \LUT[71][4] ,
         \LUT[71][3] , \LUT[71][2] , \LUT[71][1] , \LUT[71][0] , \LUT[70][15] ,
         \LUT[70][14] , \LUT[70][13] , \LUT[70][12] , \LUT[70][11] ,
         \LUT[70][10] , \LUT[70][9] , \LUT[70][8] , \LUT[70][7] , \LUT[70][6] ,
         \LUT[70][5] , \LUT[70][4] , \LUT[70][3] , \LUT[70][2] , \LUT[70][1] ,
         \LUT[70][0] , \LUT[69][15] , \LUT[69][14] , \LUT[69][13] ,
         \LUT[69][12] , \LUT[69][11] , \LUT[69][10] , \LUT[69][9] ,
         \LUT[69][8] , \LUT[69][7] , \LUT[69][6] , \LUT[69][5] , \LUT[69][4] ,
         \LUT[69][3] , \LUT[69][2] , \LUT[69][1] , \LUT[69][0] , \LUT[68][15] ,
         \LUT[68][14] , \LUT[68][13] , \LUT[68][12] , \LUT[68][11] ,
         \LUT[68][10] , \LUT[68][9] , \LUT[68][8] , \LUT[68][7] , \LUT[68][6] ,
         \LUT[68][5] , \LUT[68][4] , \LUT[68][3] , \LUT[68][2] , \LUT[68][1] ,
         \LUT[68][0] , \LUT[67][15] , \LUT[67][14] , \LUT[67][13] ,
         \LUT[67][12] , \LUT[67][11] , \LUT[67][10] , \LUT[67][9] ,
         \LUT[67][8] , \LUT[67][7] , \LUT[67][6] , \LUT[67][5] , \LUT[67][4] ,
         \LUT[67][3] , \LUT[67][2] , \LUT[67][1] , \LUT[67][0] , \LUT[66][15] ,
         \LUT[66][14] , \LUT[66][13] , \LUT[66][12] , \LUT[66][11] ,
         \LUT[66][10] , \LUT[66][9] , \LUT[66][8] , \LUT[66][7] , \LUT[66][6] ,
         \LUT[66][5] , \LUT[66][4] , \LUT[66][3] , \LUT[66][2] , \LUT[66][1] ,
         \LUT[66][0] , \LUT[65][15] , \LUT[65][14] , \LUT[65][13] ,
         \LUT[65][12] , \LUT[65][11] , \LUT[65][10] , \LUT[65][9] ,
         \LUT[65][8] , \LUT[65][7] , \LUT[65][6] , \LUT[65][5] , \LUT[65][4] ,
         \LUT[65][3] , \LUT[65][2] , \LUT[65][1] , \LUT[65][0] , \LUT[64][15] ,
         \LUT[64][14] , \LUT[64][13] , \LUT[64][12] , \LUT[64][11] ,
         \LUT[64][10] , \LUT[64][9] , \LUT[64][8] , \LUT[64][7] , \LUT[64][6] ,
         \LUT[64][5] , \LUT[64][4] , \LUT[64][3] , \LUT[64][2] , \LUT[64][1] ,
         \LUT[64][0] , \LUT[63][15] , \LUT[63][14] , \LUT[63][13] ,
         \LUT[63][12] , \LUT[63][11] , \LUT[63][10] , \LUT[63][9] ,
         \LUT[63][8] , \LUT[63][7] , \LUT[63][6] , \LUT[63][5] , \LUT[63][4] ,
         \LUT[63][3] , \LUT[63][2] , \LUT[63][1] , \LUT[63][0] , \LUT[62][15] ,
         \LUT[62][14] , \LUT[62][13] , \LUT[62][12] , \LUT[62][11] ,
         \LUT[62][10] , \LUT[62][9] , \LUT[62][8] , \LUT[62][7] , \LUT[62][6] ,
         \LUT[62][5] , \LUT[62][4] , \LUT[62][3] , \LUT[62][2] , \LUT[62][1] ,
         \LUT[62][0] , \LUT[61][15] , \LUT[61][14] , \LUT[61][13] ,
         \LUT[61][12] , \LUT[61][11] , \LUT[61][10] , \LUT[61][9] ,
         \LUT[61][8] , \LUT[61][7] , \LUT[61][6] , \LUT[61][5] , \LUT[61][4] ,
         \LUT[61][3] , \LUT[61][2] , \LUT[61][1] , \LUT[61][0] , \LUT[60][15] ,
         \LUT[60][14] , \LUT[60][13] , \LUT[60][12] , \LUT[60][11] ,
         \LUT[60][10] , \LUT[60][9] , \LUT[60][8] , \LUT[60][7] , \LUT[60][6] ,
         \LUT[60][5] , \LUT[60][4] , \LUT[60][3] , \LUT[60][2] , \LUT[60][1] ,
         \LUT[60][0] , \LUT[59][15] , \LUT[59][14] , \LUT[59][13] ,
         \LUT[59][12] , \LUT[59][11] , \LUT[59][10] , \LUT[59][9] ,
         \LUT[59][8] , \LUT[59][7] , \LUT[59][6] , \LUT[59][5] , \LUT[59][4] ,
         \LUT[59][3] , \LUT[59][2] , \LUT[59][1] , \LUT[59][0] , \LUT[58][15] ,
         \LUT[58][14] , \LUT[58][13] , \LUT[58][12] , \LUT[58][11] ,
         \LUT[58][10] , \LUT[58][9] , \LUT[58][8] , \LUT[58][7] , \LUT[58][6] ,
         \LUT[58][5] , \LUT[58][4] , \LUT[58][3] , \LUT[58][2] , \LUT[58][1] ,
         \LUT[58][0] , \LUT[57][15] , \LUT[57][14] , \LUT[57][13] ,
         \LUT[57][12] , \LUT[57][11] , \LUT[57][10] , \LUT[57][9] ,
         \LUT[57][8] , \LUT[57][7] , \LUT[57][6] , \LUT[57][5] , \LUT[57][4] ,
         \LUT[57][3] , \LUT[57][2] , \LUT[57][1] , \LUT[57][0] ,
         \LUT[119][15] , \LUT[119][14] , \LUT[119][13] , \LUT[119][12] ,
         \LUT[119][11] , \LUT[119][10] , \LUT[119][9] , \LUT[119][8] ,
         \LUT[119][7] , \LUT[119][6] , \LUT[119][5] , \LUT[119][4] ,
         \LUT[119][3] , \LUT[119][2] , \LUT[119][1] , \LUT[119][0] ,
         \LUT[118][15] , \LUT[118][14] , \LUT[118][13] , \LUT[118][12] ,
         \LUT[118][11] , \LUT[118][10] , \LUT[118][9] , \LUT[118][8] ,
         \LUT[118][7] , \LUT[118][6] , \LUT[118][5] , \LUT[118][4] ,
         \LUT[118][3] , \LUT[118][2] , \LUT[118][1] , \LUT[118][0] ,
         \LUT[117][15] , \LUT[117][14] , \LUT[117][13] , \LUT[117][12] ,
         \LUT[117][11] , \LUT[117][10] , \LUT[117][9] , \LUT[117][8] ,
         \LUT[117][7] , \LUT[117][6] , \LUT[117][5] , \LUT[117][4] ,
         \LUT[117][3] , \LUT[117][2] , \LUT[117][1] , \LUT[117][0] ,
         \LUT[116][15] , \LUT[116][14] , \LUT[116][13] , \LUT[116][12] ,
         \LUT[116][11] , \LUT[116][10] , \LUT[116][9] , \LUT[116][8] ,
         \LUT[116][7] , \LUT[116][6] , \LUT[116][5] , \LUT[116][4] ,
         \LUT[116][3] , \LUT[116][2] , \LUT[116][1] , \LUT[116][0] ,
         \LUT[115][15] , \LUT[115][14] , \LUT[115][13] , \LUT[115][12] ,
         \LUT[115][11] , \LUT[115][10] , \LUT[115][9] , \LUT[115][8] ,
         \LUT[115][7] , \LUT[115][6] , \LUT[115][5] , \LUT[115][4] ,
         \LUT[115][3] , \LUT[115][2] , \LUT[115][1] , \LUT[115][0] ,
         \LUT[114][15] , \LUT[114][14] , \LUT[114][13] , \LUT[114][12] ,
         \LUT[114][11] , \LUT[114][10] , \LUT[114][9] , \LUT[114][8] ,
         \LUT[114][7] , \LUT[114][6] , \LUT[114][5] , \LUT[114][4] ,
         \LUT[114][3] , \LUT[114][2] , \LUT[114][1] , \LUT[114][0] ,
         \LUT[113][15] , \LUT[113][14] , \LUT[113][13] , \LUT[113][12] ,
         \LUT[113][11] , \LUT[113][10] , \LUT[113][9] , \LUT[113][8] ,
         \LUT[113][7] , \LUT[113][6] , \LUT[113][5] , \LUT[113][4] ,
         \LUT[113][3] , \LUT[113][2] , \LUT[113][1] , \LUT[113][0] ,
         \LUT[112][15] , \LUT[112][14] , \LUT[112][13] , \LUT[112][12] ,
         \LUT[112][11] , \LUT[112][10] , \LUT[112][9] , \LUT[112][8] ,
         \LUT[112][7] , \LUT[112][6] , \LUT[112][5] , \LUT[112][4] ,
         \LUT[112][3] , \LUT[112][2] , \LUT[112][1] , \LUT[112][0] ,
         \LUT[111][15] , \LUT[111][14] , \LUT[111][13] , \LUT[111][12] ,
         \LUT[111][11] , \LUT[111][10] , \LUT[111][9] , \LUT[111][8] ,
         \LUT[111][7] , \LUT[111][6] , \LUT[111][5] , \LUT[111][4] ,
         \LUT[111][3] , \LUT[111][2] , \LUT[111][1] , \LUT[111][0] ,
         \LUT[110][15] , \LUT[110][14] , \LUT[110][13] , \LUT[110][12] ,
         \LUT[110][11] , \LUT[110][10] , \LUT[110][9] , \LUT[110][8] ,
         \LUT[110][7] , \LUT[110][6] , \LUT[110][5] , \LUT[110][4] ,
         \LUT[110][3] , \LUT[110][2] , \LUT[110][1] , \LUT[110][0] ,
         \LUT[109][15] , \LUT[109][14] , \LUT[109][13] , \LUT[109][12] ,
         \LUT[109][11] , \LUT[109][10] , \LUT[109][9] , \LUT[109][8] ,
         \LUT[109][7] , \LUT[109][6] , \LUT[109][5] , \LUT[109][4] ,
         \LUT[109][3] , \LUT[109][2] , \LUT[109][1] , \LUT[109][0] ,
         \LUT[108][15] , \LUT[108][14] , \LUT[108][13] , \LUT[108][12] ,
         \LUT[108][11] , \LUT[108][10] , \LUT[108][9] , \LUT[108][8] ,
         \LUT[108][7] , \LUT[108][6] , \LUT[108][5] , \LUT[108][4] ,
         \LUT[108][3] , \LUT[108][2] , \LUT[108][1] , \LUT[108][0] ,
         \LUT[107][15] , \LUT[107][14] , \LUT[107][13] , \LUT[107][12] ,
         \LUT[107][11] , \LUT[107][10] , \LUT[107][9] , \LUT[107][8] ,
         \LUT[107][7] , \LUT[107][6] , \LUT[107][5] , \LUT[107][4] ,
         \LUT[107][3] , \LUT[107][2] , \LUT[107][1] , \LUT[107][0] ,
         \LUT[106][15] , \LUT[106][14] , \LUT[106][13] , \LUT[106][12] ,
         \LUT[106][11] , \LUT[106][10] , \LUT[106][9] , \LUT[106][8] ,
         \LUT[106][7] , \LUT[106][6] , \LUT[106][5] , \LUT[106][4] ,
         \LUT[106][3] , \LUT[106][2] , \LUT[106][1] , \LUT[106][0] ,
         \LUT[105][15] , \LUT[105][14] , \LUT[105][13] , \LUT[105][12] ,
         \LUT[105][11] , \LUT[105][10] , \LUT[105][9] , \LUT[105][8] ,
         \LUT[105][7] , \LUT[105][6] , \LUT[105][5] , \LUT[105][4] ,
         \LUT[105][3] , \LUT[105][2] , \LUT[105][1] , \LUT[105][0] ,
         \LUT[104][15] , \LUT[104][14] , \LUT[104][13] , \LUT[104][12] ,
         \LUT[104][11] , \LUT[104][10] , \LUT[104][9] , \LUT[104][8] ,
         \LUT[104][7] , \LUT[104][6] , \LUT[104][5] , \LUT[104][4] ,
         \LUT[104][3] , \LUT[104][2] , \LUT[104][1] , \LUT[104][0] ,
         \LUT[103][15] , \LUT[103][14] , \LUT[103][13] , \LUT[103][12] ,
         \LUT[103][11] , \LUT[103][10] , \LUT[103][9] , \LUT[103][8] ,
         \LUT[103][7] , \LUT[103][6] , \LUT[103][5] , \LUT[103][4] ,
         \LUT[103][3] , \LUT[103][2] , \LUT[103][1] , \LUT[103][0] ,
         \LUT[102][15] , \LUT[102][14] , \LUT[102][13] , \LUT[102][12] ,
         \LUT[102][11] , \LUT[102][10] , \LUT[102][9] , \LUT[102][8] ,
         \LUT[102][7] , \LUT[102][6] , \LUT[102][5] , \LUT[102][4] ,
         \LUT[102][3] , \LUT[102][2] , \LUT[102][1] , \LUT[102][0] ,
         \LUT[101][15] , \LUT[101][14] , \LUT[101][13] , \LUT[101][12] ,
         \LUT[101][11] , \LUT[101][10] , \LUT[101][9] , \LUT[101][8] ,
         \LUT[101][7] , \LUT[101][6] , \LUT[101][5] , \LUT[101][4] ,
         \LUT[101][3] , \LUT[101][2] , \LUT[101][1] , \LUT[101][0] ,
         \LUT[100][15] , \LUT[100][14] , \LUT[100][13] , \LUT[100][12] ,
         \LUT[100][11] , \LUT[100][10] , \LUT[100][9] , \LUT[100][8] ,
         \LUT[100][7] , \LUT[100][6] , \LUT[100][5] , \LUT[100][4] ,
         \LUT[100][3] , \LUT[100][2] , \LUT[100][1] , \LUT[100][0] ,
         \LUT[99][15] , \LUT[99][14] , \LUT[99][13] , \LUT[99][12] ,
         \LUT[99][11] , \LUT[99][10] , \LUT[99][9] , \LUT[99][8] ,
         \LUT[99][7] , \LUT[99][6] , \LUT[99][5] , \LUT[99][4] , \LUT[99][3] ,
         \LUT[99][2] , \LUT[99][1] , \LUT[99][0] , \LUT[98][15] ,
         \LUT[98][14] , \LUT[98][13] , \LUT[98][12] , \LUT[98][11] ,
         \LUT[98][10] , \LUT[98][9] , \LUT[98][8] , \LUT[98][7] , \LUT[98][6] ,
         \LUT[98][5] , \LUT[98][4] , \LUT[98][3] , \LUT[98][2] , \LUT[98][1] ,
         \LUT[98][0] , \LUT[97][15] , \LUT[97][14] , \LUT[97][13] ,
         \LUT[97][12] , \LUT[97][11] , \LUT[97][10] , \LUT[97][9] ,
         \LUT[97][8] , \LUT[97][7] , \LUT[97][6] , \LUT[97][5] , \LUT[97][4] ,
         \LUT[97][3] , \LUT[97][2] , \LUT[97][1] , \LUT[97][0] , \LUT[96][15] ,
         \LUT[96][14] , \LUT[96][13] , \LUT[96][12] , \LUT[96][11] ,
         \LUT[96][10] , \LUT[96][9] , \LUT[96][8] , \LUT[96][7] , \LUT[96][6] ,
         \LUT[96][5] , \LUT[96][4] , \LUT[96][3] , \LUT[96][2] , \LUT[96][1] ,
         \LUT[96][0] , \LUT[95][15] , \LUT[95][14] , \LUT[95][13] ,
         \LUT[95][12] , \LUT[95][11] , \LUT[95][10] , \LUT[95][9] ,
         \LUT[95][8] , \LUT[95][7] , \LUT[95][6] , \LUT[95][5] , \LUT[95][4] ,
         \LUT[95][3] , \LUT[95][2] , \LUT[95][1] , \LUT[95][0] , \LUT[94][15] ,
         \LUT[94][14] , \LUT[94][13] , \LUT[94][12] , \LUT[94][11] ,
         \LUT[94][10] , \LUT[94][9] , \LUT[94][8] , \LUT[94][7] , \LUT[94][6] ,
         \LUT[94][5] , \LUT[94][4] , \LUT[94][3] , \LUT[94][2] , \LUT[94][1] ,
         \LUT[94][0] , \LUT[93][15] , \LUT[93][14] , \LUT[93][13] ,
         \LUT[93][12] , \LUT[93][11] , \LUT[93][10] , \LUT[93][9] ,
         \LUT[93][8] , \LUT[93][7] , \LUT[93][6] , \LUT[93][5] , \LUT[93][4] ,
         \LUT[93][3] , \LUT[93][2] , \LUT[93][1] , \LUT[93][0] , \LUT[92][15] ,
         \LUT[92][14] , \LUT[92][13] , \LUT[92][12] , \LUT[92][11] ,
         \LUT[92][10] , \LUT[92][9] , \LUT[92][8] , \LUT[92][7] , \LUT[92][6] ,
         \LUT[92][5] , \LUT[92][4] , \LUT[92][3] , \LUT[92][2] , \LUT[92][1] ,
         \LUT[92][0] , \LUT[91][15] , \LUT[91][14] , \LUT[91][13] ,
         \LUT[91][12] , \LUT[91][11] , \LUT[91][10] , \LUT[91][9] ,
         \LUT[91][8] , \LUT[91][7] , \LUT[91][6] , \LUT[91][5] , \LUT[91][4] ,
         \LUT[91][3] , \LUT[91][2] , \LUT[91][1] , \LUT[91][0] , \LUT[90][15] ,
         \LUT[90][14] , \LUT[90][13] , \LUT[90][12] , \LUT[90][11] ,
         \LUT[90][10] , \LUT[90][9] , \LUT[90][8] , \LUT[90][7] , \LUT[90][6] ,
         \LUT[90][5] , \LUT[90][4] , \LUT[90][3] , \LUT[90][2] , \LUT[90][1] ,
         \LUT[90][0] , \LUT[89][15] , \LUT[89][14] , \LUT[89][13] ,
         \LUT[89][12] , \LUT[89][11] , \LUT[89][10] , \LUT[89][9] ,
         \LUT[89][8] , \LUT[89][7] , \LUT[89][6] , \LUT[89][5] , \LUT[89][4] ,
         \LUT[89][3] , \LUT[89][2] , \LUT[89][1] , \LUT[89][0] , n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,
         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
         n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,
         n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
         n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,
         n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
         n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
         n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
         n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
         n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,
         n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
         n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
         n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770,
         n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778,
         n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,
         n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794,
         n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802,
         n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810,
         n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818,
         n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,
         n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834,
         n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842,
         n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850,
         n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,
         n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,
         n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874,
         n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882,
         n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890,
         n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898,
         n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906,
         n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914,
         n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922,
         n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930,
         n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938,
         n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,
         n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954,
         n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962,
         n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970,
         n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978,
         n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986,
         n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994,
         n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,
         n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010,
         n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
         n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
         n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034,
         n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
         n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,
         n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058,
         n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,
         n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
         n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
         n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
         n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
         n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106,
         n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114,
         n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,
         n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130,
         n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
         n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,
         n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154,
         n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
         n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170,
         n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178,
         n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186,
         n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194,
         n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202,
         n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
         n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218,
         n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226,
         n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
         n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,
         n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250,
         n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258,
         n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266,
         n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274,
         n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,
         n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,
         n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298,
         n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
         n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314,
         n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322,
         n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330,
         n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
         n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346,
         n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,
         n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
         n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370,
         n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
         n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,
         n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394,
         n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,
         n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
         n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
         n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
         n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
         n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,
         n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
         n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458,
         n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466,
         n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
         n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
         n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
         n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
         n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
         n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538,
         n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,
         n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
         n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562,
         n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
         n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
         n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
         n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
         n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602,
         n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610,
         n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,
         n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,
         n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634,
         n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,
         n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,
         n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658,
         n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
         n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674,
         n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682,
         n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690,
         n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
         n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706,
         n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714,
         n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722,
         n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730,
         n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
         n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746,
         n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754,
         n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762,
         n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770,
         n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778,
         n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786,
         n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,
         n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802,
         n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
         n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818,
         n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826,
         n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834,
         n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842,
         n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850,
         n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,
         n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866,
         n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874,
         n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
         n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890,
         n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898,
         n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906,
         n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914,
         n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922,
         n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,
         n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938,
         n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946,
         n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
         n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962,
         n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970,
         n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978,
         n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,
         n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,
         n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,
         n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,
         n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018,
         n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
         n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,
         n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042,
         n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050,
         n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058,
         n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
         n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074,
         n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,
         n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,
         n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
         n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106,
         n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114,
         n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122,
         n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,
         n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
         n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194,
         n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
         n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
         n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218,
         n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
         n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,
         n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
         n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250,
         n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258,
         n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266,
         n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
         n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,
         n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290,
         n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
         n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306,
         n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314,
         n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322,
         n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330,
         n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338,
         n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,
         n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
         n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362,
         n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
         n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378,
         n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386,
         n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394,
         n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402,
         n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410,
         n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,
         n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426,
         n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434,
         n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
         n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450,
         n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458,
         n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466,
         n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474,
         n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482,
         n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490,
         n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498,
         n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506,
         n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514,
         n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522,
         n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,
         n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538,
         n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546,
         n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554,
         n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,
         n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570,
         n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578,
         n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586,
         n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594,
         n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602,
         n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610,
         n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618,
         n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626,
         n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634,
         n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642,
         n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650,
         n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658,
         n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666,
         n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674,
         n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682,
         n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690,
         n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698,
         n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706,
         n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714,
         n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722,
         n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730,
         n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738,
         n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746,
         n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754,
         n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762,
         n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770,
         n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778,
         n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786,
         n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794,
         n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802,
         n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810,
         n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818,
         n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826,
         n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834,
         n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842,
         n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850,
         n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858,
         n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866,
         n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874,
         n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882,
         n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890,
         n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898,
         n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906,
         n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914,
         n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922,
         n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930,
         n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938,
         n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946,
         n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954,
         n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962,
         n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970,
         n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978,
         n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986,
         n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994,
         n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002,
         n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010,
         n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018,
         n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026,
         n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034,
         n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042,
         n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050,
         n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058,
         n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066,
         n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074,
         n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082,
         n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090,
         n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098,
         n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106,
         n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114,
         n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122,
         n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130,
         n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138,
         n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146,
         n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154,
         n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162,
         n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170,
         n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178,
         n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186,
         n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194,
         n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202,
         n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210,
         n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218,
         n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226,
         n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234,
         n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242,
         n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250,
         n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258,
         n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266,
         n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274,
         n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282,
         n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290,
         n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298,
         n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306,
         n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314,
         n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322,
         n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330,
         n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338,
         n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346,
         n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354,
         n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362,
         n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370,
         n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378,
         n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386,
         n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394,
         n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402,
         n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410,
         n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418,
         n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426,
         n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434,
         n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442,
         n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450,
         n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458,
         n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466,
         n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474,
         n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482,
         n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490,
         n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498,
         n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506,
         n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514,
         n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522,
         n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530,
         n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538,
         n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546,
         n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554,
         n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562,
         n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570,
         n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578,
         n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586,
         n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594,
         n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602,
         n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610,
         n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618,
         n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626,
         n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634,
         n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642,
         n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650,
         n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658,
         n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666,
         n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674,
         n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682,
         n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690,
         n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698,
         n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706,
         n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714,
         n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722,
         n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730,
         n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738,
         n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746,
         n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754,
         n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762,
         n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770,
         n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778,
         n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786,
         n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794,
         n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802,
         n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810,
         n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818,
         n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826,
         n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834,
         n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842,
         n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850,
         n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858,
         n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866,
         n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874,
         n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882,
         n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890,
         n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898,
         n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906,
         n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914,
         n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922,
         n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930,
         n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938,
         n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946,
         n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954,
         n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962,
         n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970,
         n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978,
         n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986,
         n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994,
         n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002,
         n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010,
         n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018,
         n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026,
         n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034,
         n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042,
         n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050,
         n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058,
         n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066,
         n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
         n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082,
         n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090,
         n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098,
         n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106,
         n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114,
         n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122,
         n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130,
         n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138,
         n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146,
         n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154,
         n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162,
         n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170,
         n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178,
         n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186,
         n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194,
         n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202,
         n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210,
         n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218,
         n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226,
         n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234,
         n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242,
         n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250,
         n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258,
         n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266,
         n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274,
         n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282,
         n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290,
         n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298,
         n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306,
         n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314,
         n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322,
         n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330,
         n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338,
         n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346,
         n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354,
         n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362,
         n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370,
         n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378,
         n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386,
         n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394,
         n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402,
         n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410,
         n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418,
         n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426,
         n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434,
         n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442,
         n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450,
         n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458,
         n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466,
         n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474,
         n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482,
         n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490,
         n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498,
         n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506,
         n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514,
         n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522,
         n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530,
         n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538,
         n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546,
         n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554,
         n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562,
         n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570,
         n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578,
         n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586,
         n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594,
         n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602,
         n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610,
         n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618,
         n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626,
         n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634,
         n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642,
         n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650,
         n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658,
         n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666,
         n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674,
         n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682,
         n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690,
         n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698,
         n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706,
         n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714,
         n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
         n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730,
         n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738,
         n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746,
         n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754,
         n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762,
         n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770,
         n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778,
         n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786,
         n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794,
         n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802,
         n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810,
         n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818,
         n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826,
         n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834,
         n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842,
         n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850,
         n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858,
         n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866,
         n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874,
         n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882,
         n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890,
         n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898,
         n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906,
         n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914,
         n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922,
         n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930,
         n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
         n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946,
         n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954,
         n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962,
         n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970,
         n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978,
         n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986,
         n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994,
         n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002,
         n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010,
         n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018,
         n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026,
         n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034,
         n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042,
         n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050,
         n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058,
         n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066,
         n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074,
         n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082,
         n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090,
         n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098,
         n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106,
         n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114,
         n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122,
         n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130,
         n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138,
         n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146,
         n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154,
         n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162,
         n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170,
         n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178,
         n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186,
         n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194,
         n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202,
         n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210,
         n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218,
         n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226,
         n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234,
         n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242,
         n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250,
         n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258,
         n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266,
         n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274,
         n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282,
         n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290,
         n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298,
         n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306,
         n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314,
         n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322,
         n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330,
         n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338,
         n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346,
         n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354,
         n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362,
         n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370,
         n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378,
         n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386,
         n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394,
         n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402,
         n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410,
         n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418,
         n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426,
         n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434,
         n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442,
         n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450,
         n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458,
         n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466,
         n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474,
         n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21482,
         n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490,
         n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498,
         n21499, n21500, n21501, n21502, n21503, n21504, n21505, n21506,
         n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514,
         n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522,
         n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530,
         n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538,
         n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546,
         n21547, n21548, n21549, n21550, n21551, n21552, n21553, n21554,
         n21555, n21556, n21557, n21558, n21559, n21560, n21561, n21562,
         n21563, n21564, n21565, n21566, n21567, n21568, n21569, n21570,
         n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578,
         n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586,
         n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594,
         n21595, n21596, n21597, n21598, n21599, n21600, n21601, n21602,
         n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610,
         n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21618,
         n21619, n21620, n21621, n21622, n21623, n21624, n21625, n21626,
         n21627, n21628, n21629, n21630, n21631, n21632, n21633, n21634,
         n21635, n21636, n21637, n21638, n21639, n21640, n21641, n21642,
         n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650,
         n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658,
         n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666,
         n21667, n21668, n21669, n21670, n21671, n21672, n21673, n21674,
         n21675, n21676, n21677, n21678, n21679, n21680, n21681, n21682,
         n21683, n21684, n21685, n21686, n21687, n21688, n21689, n21690,
         n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698,
         n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706,
         n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714,
         n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722,
         n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730,
         n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738,
         n21739, n21740, n21741, n21742, n21743, n21744, n21745, n21746,
         n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754,
         n21755, n21756, n21757, n21758, n21759, n21760, n21761, n21762,
         n21763, n21764, n21765, n21766, n21767, n21768, n21769, n21770,
         n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778,
         n21779, n21780, n21781, n21782, n21783, n21784, n21785, n21786,
         n21787, n21788, n21789, n21790, n21791, n21792, n21793, n21794,
         n21795, n21796, n21797, n21798, n21799, n21800, n21801, n21802,
         n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810,
         n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818,
         n21819, n21820, n21821, n21822, n21823, n21824, n21825, n21826,
         n21827, n21828, n21829, n21830, n21831, n21832, n21833, n21834,
         n21835, n21836, n21837, n21838, n21839, n21840, n21841, n21842,
         n21843, n21844, n21845, n21846, n21847, n21848, n21849, n21850,
         n21851, n21852, n21853, n21854, n21855, n21856, n21857, n21858,
         n21859, n21860, n21861, n21862, n21863, n21864, n21865, n21866,
         n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874,
         n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882,
         n21883, n21884, n21885, n21886, n21887, n21888, n21889, n21890,
         n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898,
         n21899, n21900, n21901, n21902, n21903, n21904, n21905, n21906,
         n21907, n21908, n21909, n21910, n21911, n21912, n21913, n21914,
         n21915, n21916, n21917, n21918, n21919, n21920, n21921, n21922,
         n21923, n21924, n21925, n21926, n21927, n21928, n21929, n21930,
         n21931, n21932, n21933, n21934, n21935, n21936, n21937, n21938,
         n21939, n21940, n21941, n21942, n21943, n21944, n21945, n21946,
         n21947, n21948, n21949, n21950, n21951, n21952, n21953, n21954,
         n21955, n21956, n21957, n21958, n21959, n21960, n21961, n21962,
         n21963, n21964, n21965, n21966, n21967, n21968, n21969, n21970,
         n21971, n21972, n21973, n21974, n21975, n21976, n21977, n21978,
         n21979, n21980, n21981, n21982, n21983, n21984, n21985, n21986,
         n21987, n21988, n21989, n21990, n21991, n21992, n21993, n21994,
         n21995, n21996, n21997, n21998, n21999, n22000, n22001, n22002,
         n22003, n22004, n22005, n22006, n22007, n22008, n22009, n22010,
         n22011, n22012, n22013, n22014, n22015, n22016, n22017, n22018,
         n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026,
         n22027, n22028, n22029, n22030, n22031, n22032, n22033, n22034,
         n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042,
         n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050,
         n22051, n22052, n22053, n22054, n22055, n22056, n22057, n22058,
         n22059, n22060, n22061, n22062, n22063, n22064, n22065, n22066,
         n22067, n22068, n22069, n22070, n22071, n22072, n22073, n22074,
         n22075, n22076, n22077, n22078, n22079, n22080, n22081, n22082,
         n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090,
         n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098,
         n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106,
         n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114,
         n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122,
         n22123, n22124, n22125, n22126, n22127, n22128, n22129, n22130,
         n22131, n22132, n22133, n22134, n22135, n22136, n22137, n22138,
         n22139, n22140, n22141, n22142, n22143, n22144, n22145, n22146,
         n22147, n22148, n22149, n22150, n22151, n22152, n22153, n22154,
         n22155, n22156, n22157, n22158, n22159, n22160, n22161, n22162,
         n22163, n22164, n22165, n22166, n22167, n22168, n22169, n22170,
         n22171, n22172, n22173, n22174, n22175, n22176, n22177, n22178,
         n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186,
         n22187, n22188, n22189, n22190, n22191, n22192, n22193, n22194,
         n22195, n22196, n22197, n22198, n22199, n22200, n22201, n22202,
         n22203, n22204, n22205, n22206, n22207, n22208, n22209, n22210,
         n22211, n22212, n22213, n22214, n22215, n22216, n22217, n22218,
         n22219, n22220, n22221, n22222, n22223, n22224, n22225, n22226,
         n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234,
         n22235, n22236, n22237, n22238, n22239, n22240, n22241, n22242,
         n22243, n22244, n22245, n22246, n22247, n22248, n22249, n22250,
         n22251, n22252, n22253, n22254, n22255, n22256, n22257, n22258,
         n22259, n22260, n22261, n22262, n22263, n22264, n22265, n22266,
         n22267, n22268, n22269, n22270, n22271, n22272, n22273, n22274,
         n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282,
         n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22290,
         n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298,
         n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306,
         n22307, n22308, n22309, n22310, n22311, n22312, n22313, n22314,
         n22315, n22316, n22317, n22318, n22319, n22320, n22321, n22322,
         n22323, n22324, n22325, n22326, n22327, n22328, n22329, n22330,
         n22331, n22332, n22333, n22334, n22335, n22336, n22337, n22338,
         n22339, n22340, n22341, n22342, n22343, n22344, n22345, n22346,
         n22347, n22348, n22349, n22350, n22351, n22352, n22353, n22354,
         n22355, n22356, n22357, n22358, n22359, n22360, n22361, n22362,
         n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370,
         n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378,
         n22379, n22380, n22381, n22382, n22383, n22384, n22385, n22386,
         n22387, n22388, n22389, n22390, n22391, n22392, n22393, n22394,
         n22395, n22396, n22397, n22398, n22399, n22400, n22401, n22402,
         n22403, n22404, n22405, n22406, n22407, n22408, n22409, n22410,
         n22411, n22412, n22413, n22414, n22415, n22416, n22417, n22418,
         n22419, n22420, n22421, n22422, n22423, n22424, n22425, n22426,
         n22427, n22428, n22429, n22430, n22431, n22432, n22433, n22434,
         n22435, n22436, n22437, n22438, n22439, n22440, n22441, n22442,
         n22443, n22444, n22445, n22446, n22447, n22448, n22449, n22450,
         n22451, n22452, n22453, n22454, n22455, n22456, n22457, n22458,
         n22459, n22460, n22461, n22462, n22463, n22464, n22465, n22466,
         n22467, n22468, n22469, n22470, n22471, n22472, n22473, n22474,
         n22475, n22476, n22477, n22478, n22479, n22480, n22481, n22482,
         n22483, n22484, n22485, n22486, n22487, n22488, n22489, n22490,
         n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498,
         n22499, n22500, n22501, n22502, n22503, n22504, n22505, n22506,
         n22507, n22508, n22509, n22510, n22511, n22512, n22513, n22514,
         n22515, n22516, n22517, n22518, n22519, n22520, n22521, n22522,
         n22523, n22524, n22525, n22526, n22527, n22528, n22529, n22530,
         n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538,
         n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546,
         n22547, n22548, n22549, n22550, n22551, n22552, n22553, n22554,
         n22555, n22556, n22557, n22558, n22559, n22560, n22561, n22562,
         n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570,
         n22571, n22572, n22573, n22574, n22575, n22576, n22577, n22578,
         n22579, n22580, n22581, n22582, n22583, n22584, n22585, n22586,
         n22587, n22588, n22589, n22590, n22591, n22592, n22593, n22594,
         n22595, n22596, n22597, n22598, n22599, n22600, n22601, n22602,
         n22603, n22604, n22605, n22606, n22607, n22608, n22609, n22610,
         n22611, n22612, n22613, n22614, n22615, n22616, n22617, n22618,
         n22619, n22620, n22621, n22622, n22623, n22624, n22625, n22626,
         n22627, n22628, n22629, n22630, n22631, n22632, n22633, n22634,
         n22635, n22636, n22637, n22638, n22639, n22640, n22641, n22642,
         n22643, n22644, n22645, n22646, n22647, n22648, n22649, n22650,
         n22651, n22652, n22653, n22654, n22655, n22656, n22657, n22658,
         n22659, n22660, n22661, n22662, n22663, n22664, n22665, n22666,
         n22667, n22668, n22669, n22670, n22671, n22672, n22673, n22674,
         n22675, n22676, n22677, n22678, n22679, n22680, n22681, n22682,
         n22683, n22684, n22685, n22686, n22687, n22688, n22689, n22690,
         n22691, n22692, n22693, n22694, n22695, n22696, n22697, n22698,
         n22699, n22700, n22701, n22702, n22703, n22704, n22705, n22706,
         n22707, n22708, n22709, n22710, n22711, n22712, n22713, n22714,
         n22715, n22716, n22717, n22718, n22719, n22720, n22721, n22722,
         n22723, n22724, n22725, n22726, n22727, n22728, n22729, n22730,
         n22731, n22732, n22733, n22734, n22735, n22736, n22737, n22738,
         n22739, n22740, n22741, n22742, n22743, n22744, n22745, n22746,
         n22747, n22748, n22749, n22750, n22751, n22752, n22753, n22754,
         n22755, n22756, n22757, n22758, n22759, n22760, n22761, n22762,
         n22763, n22764, n22765, n22766, n22767, n22768, n22769, n22770,
         n22771, n22772, n22773, n22774, n22775, n22776, n22777, n22778,
         n22779, n22780, n22781, n22782, n22783, n22784, n22785, n22786,
         n22787, n22788, n22789, n22790, n22791, n22792, n22793, n22794,
         n22795, n22796, n22797, n22798, n22799, n22800, n22801, n22802,
         n22803, n22804, n22805, n22806, n22807, n22808, n22809, n22810,
         n22811, n22812, n22813, n22814, n22815, n22816, n22817, n22818,
         n22819, n22820, n22821, n22822, n22823, n22824, n22825, n22826,
         n22827, n22828, n22829, n22830, n22831, n22832, n22833, n22834,
         n22835, n22836, n22837, n22838, n22839, n22840, n22841, n22842,
         n22843, n22844, n22845, n22846, n22847, n22848, n22849, n22850,
         n22851, n22852, n22853, n22854, n22855, n22856, n22857, n22858,
         n22859, n22860, n22861, n22862, n22863, n22864, n22865, n22866,
         n22867, n22868, n22869, n22870, n22871, n22872, n22873, n22874,
         n22875, n22876, n22877, n22878, n22879, n22880, n22881, n22882,
         n22883, n22884, n22885, n22886, n22887, n22888, n22889, n22890,
         n22891, n22892, n22893, n22894, n22895, n22896, n22897, n22898,
         n22899, n22900, n22901, n22902, n22903, n22904, n22905, n22906,
         n22907, n22908, n22909, n22910, n22911, n22912, n22913, n22914,
         n22915, n22916, n22917, n22918, n22919, n22920, n22921, n22922,
         n22923, n22924, n22925, n22926, n22927, n22928, n22929, n22930,
         n22931, n22932, n22933, n22934, n22935, n22936, n22937, n22938,
         n22939, n22940, n22941, n22942, n22943, n22944, n22945, n22946,
         n22947, n22948, n22949, n22950, n22951, n22952, n22953, n22954,
         n22955, n22956, n22957, n22958, n22959, n22960, n22961, n22962,
         n22963, n22964, n22965, n22966, n22967, n22968, n22969, n22970,
         n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22978,
         n22979, n22980, n22981, n22982, n22983, n22984, n22985, n22986,
         n22987, n22988, n22989, n22990, n22991, n22992, n22993, n22994,
         n22995, n22996, n22997, n22998, n22999, n23000, n23001, n23002,
         n23003, n23004, n23005, n23006, n23007, n23008, n23009, n23010,
         n23011, n23012, n23013, n23014, n23015, n23016, n23017, n23018,
         n23019, n23020, n23021, n23022, n23023, n23024, n23025, n23026,
         n23027, n23028, n23029, n23030, n23031, n23032, n23033, n23034,
         n23035, n23036, n23037, n23038, n23039, n23040, n23041, n23042,
         n23043, n23044, n23045, n23046, n23047, n23048, n23049, n23050,
         n23051, n23052, n23053, n23054, n23055, n23056, n23057, n23058,
         n23059, n23060, n23061, n23062, n23063, n23064, n23065, n23066,
         n23067, n23068, n23069, n23070, n23071, n23072, n23073, n23074,
         n23075, n23076, n23077, n23078, n23079, n23080, n23081, n23082,
         n23083, n23084, n23085, n23086, n23087, n23088, n23089, n23090,
         n23091, n23092, n23093, n23094, n23095, n23096, n23097, n23098,
         n23099, n23100, n23101, n23102, n23103, n23104, n23105, n23106,
         n23107, n23108, n23109, n23110, n23111, n23112, n23113, n23114,
         n23115, n23116, n23117, n23118, n23119, n23120, n23121, n23122,
         n23123, n23124, n23125, n23126, n23127, n23128, n23129, n23130,
         n23131, n23132, n23133, n23134, n23135, n23136, n23137, n23138,
         n23139, n23140, n23141, n23142, n23143, n23144, n23145, n23146,
         n23147, n23148, n23149, n23150, n23151, n23152, n23153, n23154,
         n23155, n23156, n23157, n23158, n23159, n23160, n23161, n23162,
         n23163, n23164, n23165, n23166, n23167, n23168, n23169, n23170,
         n23171, n23172, n23173, n23174, n23175, n23176, n23177, n23178,
         n23179, n23180, n23181, n23182, n23183, n23184, n23185, n23186,
         n23187, n23188, n23189, n23190, n23191, n23192, n23193, n23194,
         n23195, n23196, n23197, n23198, n23199, n23200, n23201, n23202,
         n23203, n23204, n23205, n23206, n23207, n23208, n23209, n23210,
         n23211, n23212, n23213, n23214, n23215, n23216, n23217, n23218,
         n23219, n23220, n23221, n23222, n23223, n23224, n23225, n23226,
         n23227, n23228, n23229, n23230, n23231, n23232, n23233, n23234,
         n23235, n23236, n23237, n23238, n23239, n23240, n23241, n23242,
         n23243, n23244, n23245, n23246, n23247, n23248, n23249, n23250,
         n23251, n23252, n23253, n23254, n23255, n23256, n23257, n23258,
         n23259, n23260, n23261, n23262, n23263, n23264, n23265, n23266,
         n23267, n23268, n23269, n23270, n23271, n23272, n23273, n23274,
         n23275, n23276, n23277, n23278, n23279, n23280, n23281, n23282,
         n23283, n23284, n23285, n23286, n23287, n23288, n23289, n23290,
         n23291, n23292, n23293, n23294, n23295, n23296, n23297, n23298,
         n23299, n23300, n23301, n23302, n23303, n23304, n23305, n23306,
         n23307, n23308, n23309, n23310, n23311, n23312, n23313, n23314,
         n23315, n23316, n23317, n23318, n23319, n23320, n23321, n23322,
         n23323, n23324, n23325, n23326, n23327, n23328, n23329, n23330,
         n23331, n23332, n23333, n23334, n23335, n23336, n23337, n23338,
         n23339, n23340, n23341, n23342, n23343, n23344, n23345, n23346,
         n23347, n23348, n23349, n23350, n23351, n23352, n23353, n23354,
         n23355, n23356, n23357, n23358, n23359, n23360, n23361, n23362,
         n23363, n23364, n23365, n23366, n23367, n23368, n23369, n23370,
         n23371, n23372, n23373, n23374, n23375, n23376, n23377, n23378,
         n23379, n23380, n23381, n23382, n23383, n23384, n23385, n23386,
         n23387, n23388, n23389, n23390, n23391, n23392, n23393, n23394,
         n23395, n23396, n23397, n23398, n23399, n23400, n23401, n23402,
         n23403, n23404, n23405, n23406, n23407, n23408, n23409, n23410,
         n23411, n23412, n23413, n23414, n23415, n23416, n23417, n23418,
         n23419, n23420, n23421, n23422, n23423, n23424, n23425, n23426,
         n23427, n23428, n23429, n23430, n23431, n23432, n23433, n23434,
         n23435, n23436, n23437, n23438, n23439, n23440, n23441, n23442,
         n23443, n23444, n23445, n23446, n23447, n23448, n23449, n23450,
         n23451, n23452, n23453, n23454, n23455, n23456, n23457, n23458,
         n23459, n23460, n23461, n23462, n23463, n23464, n23465, n23466,
         n23467, n23468, n23469, n23470, n23471, n23472, n23473, n23474,
         n23475, n23476, n23477, n23478, n23479, n23480, n23481, n23482,
         n23483, n23484, n23485, n23486, n23487, n23488, n23489, n23490,
         n23491, n23492, n23493, n23494, n23495, n23496, n23497, n23498,
         n23499, n23500, n23501, n23502, n23503, n23504, n23505, n23506,
         n23507, n23508, n23509, n23510, n23511, n23512, n23513, n23514,
         n23515, n23516, n23517, n23518, n23519, n23520, n23521, n23522,
         n23523, n23524, n23525, n23526, n23527, n23528, n23529, n23530,
         n23531, n23532, n23533, n23534, n23535, n23536, n23537, n23538,
         n23539, n23540, n23541, n23542, n23543, n23544, n23545, n23546,
         n23547, n23548, n23549, n23550, n23551, n23552, n23553, n23554,
         n23555, n23556, n23557, n23558, n23559, n23560, n23561, n23562,
         n23563, n23564, n23565, n23566, n23567, n23568, n23569, n23570,
         n23571, n23572, n23573, n23574, n23575, n23576, n23577, n23578,
         n23579, n23580, n23581, n23582, n23583, n23584, n23585, n23586,
         n23587, n23588, n23589, n23590, n23591, n23592, n23593, n23594,
         n23595, n23596, n23597, n23598, n23599, n23600, n23601, n23602,
         n23603, n23604, n23605, n23606, n23607, n23608, n23609, n23610,
         n23611, n23612, n23613, n23614, n23615, n23616, n23617, n23618,
         n23619, n23620, n23621, n23622, n23623, n23624, n23625, n23626,
         n23627, n23628, n23629, n23630, n23631, n23632, n23633, n23634,
         n23635, n23636, n23637, n23638, n23639, n23640, n23641, n23642,
         n23643, n23644, n23645, n23646, n23647, n23648, n23649, n23650,
         n23651, n23652, n23653, n23654, n23655, n23656, n23657, n23658,
         n23659, n23660, n23661, n23662, n23663, n23664, n23665, n23666,
         n23667, n23668, n23669, n23670, n23671, n23672, n23673, n23674,
         n23675, n23676, n23677, n23678, n23679, n23680, n23681, n23682,
         n23683, n23684, n23685, n23686, n23687, n23688, n23689, n23690,
         n23691, n23692, n23693, n23694, n23695, n23696, n23697, n23698,
         n23699, n23700, n23701, n23702, n23703, n23704, n23705, n23706,
         n23707, n23708, n23709, n23710, n23711, n23712, n23713, n23714,
         n23715, n23716, n23717, n23718, n23719, n23720, n23721, n23722,
         n23723, n23724, n23725, n23726, n23727, n23728, n23729, n23730,
         n23731, n23732, n23733, n23734, n23735, n23736, n23737, n23738,
         n23739, n23740, n23741, n23742, n23743, n23744, n23745, n23746,
         n23747, n23748, n23749, n23750, n23751, n23752, n23753, n23754,
         n23755, n23756, n23757, n23758, n23759, n23760, n23761, n23762,
         n23763, n23764, n23765, n23766, n23767, n23768, n23769, n23770,
         n23771, n23772, n23773, n23774, n23775, n23776, n23777, n23778,
         n23779, n23780, n23781, n23782, n23783, n23784, n23785, n23786,
         n23787, n23788, n23789, n23790, n23791, n23792, n23793, n23794,
         n23795, n23796, n23797, n23798, n23799, n23800, n23801, n23802,
         n23803, n23804, n23805, n23806, n23807, n23808, n23809, n23810,
         n23811, n23812, n23813, n23814, n23815, n23816, n23817, n23818,
         n23819, n23820, n23821, n23822, n23823, n23824, n23825, n23826,
         n23827, n23828, n23829, n23830, n23831, n23832, n23833, n23834,
         n23835, n23836, n23837, n23838, n23839, n23840, n23841, n23842,
         n23843, n23844, n23845, n23846, n23847, n23848, n23849, n23850,
         n23851, n23852, n23853, n23854, n23855, n23856, n23857, n23858,
         n23859, n23860, n23861, n23862, n23863, n23864, n23865, n23866,
         n23867, n23868, n23869, n23870, n23871, n23872, n23873, n23874,
         n23875, n23876, n23877, n23878, n23879, n23880, n23881, n23882,
         n23883, n23884, n23885, n23886, n23887, n23888, n23889, n23890,
         n23891, n23892, n23893, n23894, n23895, n23896, n23897, n23898,
         n23899, n23900, n23901, n23902, n23903, n23904, n23905, n23906,
         n23907, n23908, n23909, n23910, n23911, n23912, n23913, n23914,
         n23915, n23916, n23917, n23918, n23919, n23920, n23921, n23922,
         n23923, n23924, n23925, n23926, n23927, n23928, n23929, n23930,
         n23931, n23932, n23933, n23934, n23935, n23936, n23937, n23938,
         n23939, n23940, n23941, n23942, n23943, n23944, n23945, n23946,
         n23947, n23948, n23949, n23950, n23951, n23952, n23953, n23954,
         n23955, n23956, n23957, n23958, n23959, n23960, n23961, n23962,
         n23963, n23964, n23965, n23966, n23967, n23968, n23969, n23970,
         n23971, n23972, n23973, n23974, n23975, n23976, n23977, n23978,
         n23979, n23980, n23981, n23982, n23983, n23984, n23985, n23986,
         n23987, n23988, n23989, n23990, n23991, n23992, n23993, n23994,
         n23995, n23996, n23997, n23998, n23999, n24000, n24001, n24002,
         n24003, n24004, n24005, n24006, n24007, n24008, n24009, n24010,
         n24011, n24012, n24013, n24014, n24015, n24016, n24017, n24018,
         n24019, n24020, n24021, n24022, n24023, n24024, n24025, n24026,
         n24027, n24028, n24029, n24030, n24031, n24032, n24033, n24034,
         n24035, n24036, n24037, n24038, n24039, n24040, n24041, n24042,
         n24043, n24044, n24045, n24046, n24047, n24048, n24049, n24050,
         n24051, n24052, n24053, n24054, n24055, n24056, n24057, n24058,
         n24059, n24060, n24061, n24062, n24063, n24064, n24065, n24066,
         n24067, n24068, n24069, n24070, n24071, n24072, n24073, n24074,
         n24075, n24076, n24077, n24078, n24079, n24080, n24081, n24082,
         n24083, n24084, n24085, n24086, n24087, n24088, n24089, n24090,
         n24091, n24092, n24093, n24094, n24095, n24096, n24097, n24098,
         n24099, n24100, n24101, n24102, n24103, n24104, n24105, n24106,
         n24107, n24108, n24109, n24110, n24111, n24112, n24113, n24114,
         n24115, n24116, n24117, n24118, n24119, n24120, n24121, n24122,
         n24123, n24124, n24125, n24126, n24127, n24128, n24129, n24130,
         n24131, n24132, n24133, n24134, n24135, n24136, n24137, n24138,
         n24139, n24140, n24141, n24142, n24143, n24144, n24145, n24146,
         n24147, n24148, n24149, n24150, n24151, n24152, n24153, n24154,
         n24155, n24156, n24157, n24158, n24159, n24160, n24161, n24162,
         n24163, n24164, n24165, n24166, n24167, n24168, n24169, n24170,
         n24171, n24172, n24173, n24174, n24175, n24176, n24177, n24178,
         n24179, n24180, n24181, n24182, n24183, n24184, n24185, n24186,
         n24187, n24188, n24189, n24190, n24191, n24192, n24193, n24194,
         n24195, n24196, n24197, n24198, n24199, n24200, n24201, n24202,
         n24203, n24204, n24205, n24206, n24207, n24208, n24209, n24210,
         n24211, n24212, n24213, n24214, n24215, n24216, n24217, n24218,
         n24219, n24220, n24221, n24222, n24223, n24224, n24225, n24226,
         n24227, n24228, n24229, n24230, n24231, n24232, n24233, n24234,
         n24235, n24236, n24237, n24238, n24239, n24240, n24241, n24242,
         n24243, n24244, n24245, n24246, n24247, n24248, n24249, n24250,
         n24251, n24252, n24253, n24254, n24255, n24256, n24257, n24258,
         n24259, n24260, n24261, n24262, n24263, n24264, n24265, n24266,
         n24267, n24268, n24269, n24270, n24271, n24272, n24273, n24274,
         n24275, n24276, n24277, n24278, n24279, n24280, n24281, n24282,
         n24283, n24284, n24285, n24286, n24287, n24288, n24289, n24290,
         n24291, n24292, n24293, n24294, n24295, n24296, n24297, n24298,
         n24299, n24300, n24301, n24302, n24303, n24304, n24305, n24306,
         n24307, n24308, n24309, n24310, n24311, n24312, n24313, n24314,
         n24315, n24316, n24317, n24318, n24319, n24320, n24321, n24322,
         n24323, n24324, n24325, n24326, n24327, n24328, n24329, n24330,
         n24331, n24332, n24333, n24334, n24335, n24336, n24337, n24338,
         n24339, n24340, n24341, n24342, n24343, n24344, n24345, n24346,
         n24347, n24348, n24349, n24350, n24351, n24352, n24353, n24354,
         n24355, n24356, n24357, n24358, n24359, n24360, n24361, n24362,
         n24363, n24364, n24365, n24366, n24367, n24368, n24369, n24370,
         n24371, n24372, n24373, n24374, n24375, n24376, n24377, n24378,
         n24379, n24380, n24381, n24382, n24383, n24384, n24385, n24386,
         n24387, n24388, n24389, n24390, n24391, n24392, n24393, n24394,
         n24395, n24396, n24397, n24398, n24399, n24400, n24401, n24402,
         n24403, n24404, n24405, n24406, n24407, n24408, n24409, n24410,
         n24411, n24412, n24413, n24414, n24415, n24416, n24417, n24418,
         n24419, n24420, n24421, n24422, n24423, n24424, n24425, n24426,
         n24427, n24428, n24429, n24430, n24431, n24432, n24433, n24434,
         n24435, n24436, n24437, n24438, n24439, n24440, n24441, n24442,
         n24443, n24444, n24445, n24446, n24447, n24448, n24449, n24450,
         n24451, n24452, n24453, n24454, n24455, n24456, n24457, n24458,
         n24459, n24460, n24461, n24462, n24463, n24464, n24465, n24466,
         n24467, n24468, n24469, n24470, n24471, n24472, n24473, n24474,
         n24475, n24476, n24477, n24478, n24479, n24480, n24481, n24482,
         n24483, n24484, n24485, n24486, n24487, n24488, n24489, n24490,
         n24491, n24492, n24493, n24494, n24495, n24496, n24497, n24498,
         n24499, n24500, n24501, n24502, n24503, n24504, n24505, n24506,
         n24507, n24508, n24509, n24510, n24511, n24512, n24513, n24514,
         n24515, n24516, n24517, n24518, n24519, n24520, n24521, n24522,
         n24523, n24524, n24525, n24526, n24527, n24528, n24529, n24530,
         n24531, n24532, n24533, n24534, n24535, n24536, n24537, n24538,
         n24539, n24540, n24541, n24542, n24543, n24544, n24545, n24546,
         n24547, n24548, n24549, n24550, n24551, n24552, n24553, n24554,
         n24555, n24556, n24557, n24558, n24559, n24560, n24561, n24562,
         n24563, n24564, n24565, n24566, n24567, n24568, n24569, n24570,
         n24571, n24572, n24573, n24574, n24575, n24576, n24577, n24578,
         n24579, n24580, n24581, n24582, n24583, n24584, n24585, n24586,
         n24587, n24588, n24589, n24590, n24591, n24592, n24593, n24594,
         n24595, n24596, n24597, n24598, n24599, n24600, n24601, n24602,
         n24603, n24604, n24605, n24606, n24607, n24608, n24609, n24610,
         n24611, n24612, n24613, n24614, n24615, n24616, n24617, n24618,
         n24619, n24620, n24621, n24622, n24623, n24624, n24625, n24626,
         n24627, n24628, n24629, n24630, n24631, n24632, n24633, n24634,
         n24635, n24636, n24637, n24638, n24639, n24640, n24641, n24642,
         n24643, n24644, n24645, n24646, n24647, n24648, n24649, n24650,
         n24651, n24652, n24653, n24654, n24655, n24656, n24657, n24658,
         n24659, n24660, n24661, n24662, n24663, n24664, n24665, n24666,
         n24667, n24668, n24669, n24670, n24671, n24672, n24673, n24674,
         n24675, n24676, n24677, n24678, n24679, n24680, n24681, n24682,
         n24683, n24684, n24685, n24686, n24687, n24688, n24689, n24690,
         n24691, n24692, n24693, n24694, n24695, n24696, n24697, n24698,
         n24699, n24700, n24701, n24702, n24703, n24704, n24705, n24706,
         n24707, n24708, n24709, n24710, n24711, n24712, n24713, n24714,
         n24715, n24716, n24717, n24718, n24719, n24720, n24721, n24722,
         n24723, n24724, n24725, n24726, n24727, n24728, n24729, n24730,
         n24731, n24732, n24733, n24734, n24735, n24736, n24737, n24738,
         n24739, n24740, n24741, n24742, n24743, n24744, n24745, n24746,
         n24747, n24748, n24749, n24750, n24751, n24752, n24753, n24754,
         n24755, n24756, n24757, n24758, n24759, n24760, n24761, n24762,
         n24763, n24764, n24765, n24766, n24767, n24768, n24769, n24770,
         n24771, n24772, n24773, n24774, n24775, n24776, n24777, n24778,
         n24779, n24780, n24781, n24782, n24783, n24784, n24785, n24786,
         n24787, n24788, n24789, n24790, n24791, n24792, n24793, n24794,
         n24795, n24796, n24797, n24798, n24799, n24800, n24801, n24802,
         n24803, n24804, n24805, n24806, n24807, n24808, n24809, n24810,
         n24811, n24812, n24813, n24814, n24815, n24816, n24817, n24818,
         n24819, n24820, n24821, n24822, n24823, n24824, n24825, n24826,
         n24827, n24828, n24829, n24830, n24831, n24832, n24833, n24834,
         n24835, n24836, n24837, n24838, n24839, n24840, n24841, n24842,
         n24843, n24844, n24845, n24846, n24847, n24848, n24849, n24850,
         n24851, n24852, n24853, n24854, n24855, n24856, n24857, n24858,
         n24859, n24860, n24861, n24862, n24863, n24864, n24865, n24866,
         n24867, n24868, n24869, n24870, n24871, n24872, n24873, n24874,
         n24875, n24876, n24877, n24878, n24879, n24880, n24881, n24882,
         n24883, n24884, n24885, n24886, n24887, n24888, n24889, n24890,
         n24891, n24892, n24893, n24894, n24895, n24896, n24897, n24898,
         n24899, n24900, n24901, n24902, n24903, n24904, n24905, n24906,
         n24907, n24908, n24909, n24910, n24911, n24912, n24913, n24914,
         n24915, n24916, n24917, n24918, n24919, n24920, n24921, n24922,
         n24923, n24924, n24925, n24926, n24927, n24928, n24929, n24930,
         n24931, n24932, n24933, n24934, n24935, n24936, n24937, n24938,
         n24939, n24940, n24941, n24942, n24943, n24944, n24945, n24946,
         n24947, n24948, n24949, n24950, n24951, n24952, n24953, n24954,
         n24955, n24956, n24957, n24958, n24959, n24960, n24961, n24962,
         n24963, n24964, n24965, n24966, n24967, n24968, n24969, n24970,
         n24971, n24972, n24973, n24974, n24975, n24976, n24977, n24978,
         n24979, n24980, n24981, n24982, n24983, n24984, n24985, n24986,
         n24987, n24988, n24989, n24990, n24991, n24992, n24993, n24994,
         n24995, n24996, n24997, n24998, n24999, n25000, n25001, n25002,
         n25003, n25004, n25005, n25006, n25007, n25008, n25009, n25010,
         n25011, n25012, n25013, n25014, n25015, n25016, n25017, n25018,
         n25019, n25020, n25021, n25022, n25023, n25024, n25025, n25026,
         n25027, n25028, n25029, n25030, n25031, n25032, n25033, n25034,
         n25035, n25036, n25037, n25038, n25039, n25040, n25041, n25042,
         n25043, n25044, n25045, n25046, n25047, n25048, n25049, n25050,
         n25051, n25052, n25053, n25054, n25055, n25056, n25057, n25058,
         n25059, n25060, n25061, n25062, n25063, n25064, n25065, n25066,
         n25067, n25068, n25069, n25070, n25071, n25072, n25073, n25074,
         n25075, n25076, n25077, n25078, n25079, n25080, n25081, n25082,
         n25083, n25084, n25085, n25086, n25087, n25088, n25089, n25090,
         n25091, n25092, n25093, n25094, n25095, n25096, n25097, n25098,
         n25099, n25100, n25101, n25102, n25103, n25104, n25105, n25106,
         n25107, n25108, n25109, n25110, n25111, n25112, n25113, n25114,
         n25115, n25116, n25117, n25118, n25119, n25120, n25121, n25122,
         n25123, n25124, n25125, n25126, n25127, n25128, n25129, n25130,
         n25131, n25132, n25133, n25134, n25135, n25136, n25137, n25138,
         n25139, n25140, n25141, n25142, n25143, n25144, n25145, n25146,
         n25147, n25148, n25149, n25150, n25151, n25152, n25153, n25154,
         n25155, n25156, n25157, n25158, n25159, n25160, n25161, n25162,
         n25163, n25164, n25165, n25166, n25167, n25168, n25169, n25170,
         n25171, n25172, n25173, n25174, n25175, n25176, n25177, n25178,
         n25179, n25180, n25181, n25182, n25183, n25184, n25185, n25186,
         n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194,
         n25195, n25196, n25197, n25198, n25199, n25200, n25201, n25202,
         n25203, n25204, n25205, n25206, n25207, n25208, n25209, n25210,
         n25211, n25212, n25213, n25214, n25215, n25216, n25217, n25218,
         n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226,
         n25227, n25228, n25229, n25230, n25231, n25232, n25233, n25234,
         n25235, n25236, n25237, n25238, n25239, n25240, n25241, n25242,
         n25243, n25244, n25245, n25246, n25247, n25248, n25249, n25250,
         n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258,
         n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266,
         n25267, n25268, n25269, n25270, n25271, n25272, n25273, n25274,
         n25275, n25276, n25277, n25278, n25279, n25280, n25281, n25282,
         n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290,
         n25291, n25292, n25293, n25294, n25295, n25296, n25297, n25298,
         n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306,
         n25307, n25308, n25309, n25310, n25311, n25312, n25313, n25314,
         n25315, n25316, n25317, n25318, n25319, n25320, n25321, n25322,
         n25323, n25324, n25325, n25326, n25327, n25328, n25329, n25330,
         n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338,
         n25339, n25340, n25341, n25342, n25343, n25344, n25345, n25346,
         n25347, n25348, n25349, n25350, n25351, n25352, n25353, n25354,
         n25355, n25356, n25357, n25358, n25359, n25360, n25361, n25362,
         n25363, n25364, n25365, n25366, n25367, n25368, n25369, n25370,
         n25371, n25372, n25373, n25374, n25375, n25376, n25377, n25378,
         n25379, n25380, n25381, n25382, n25383, n25384, n25385, n25386,
         n25387, n25388, n25389, n25390, n25391, n25392, n25393, n25394,
         n25395, n25396, n25397, n25398, n25399, n25400, n25401, n25402,
         n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410,
         n25411, n25412, n25413, n25414, n25415, n25416, n25417, n25418,
         n25419, n25420, n25421, n25422, n25423, n25424, n25425, n25426,
         n25427, n25428, n25429, n25430, n25431, n25432, n25433, n25434,
         n25435, n25436, n25437, n25438, n25439, n25440, n25441, n25442,
         n25443, n25444, n25445, n25446, n25447, n25448, n25449, n25450,
         n25451, n25452, n25453, n25454, n25455, n25456, n25457, n25458,
         n25459, n25460, n25461, n25462, n25463, n25464, n25465, n25466,
         n25467, n25468, n25469, n25470, n25471, n25472, n25473, n25474,
         n25475, n25476, n25477, n25478, n25479, n25480, n25481, n25482,
         n25483, n25484, n25485, n25486, n25487, n25488, n25489, n25490,
         n25491, n25492, n25493, n25494, n25495, n25496, n25497, n25498,
         n25499, n25500, n25501, n25502, n25503, n25504, n25505, n25506,
         n25507, n25508, n25509, n25510, n25511, n25512, n25513, n25514,
         n25515, n25516, n25517, n25518, n25519, n25520, n25521, n25522,
         n25523, n25524, n25525, n25526, n25527, n25528, n25529, n25530,
         n25531, n25532, n25533, n25534, n25535, n25536, n25537, n25538,
         n25539, n25540, n25541, n25542, n25543, n25544, n25545, n25546,
         n25547, n25548, n25549, n25550, n25551, n25552, n25553, n25554,
         n25555, n25556, n25557, n25558, n25559, n25560, n25561, n25562,
         n25563, n25564, n25565, n25566, n25567, n25568, n25569, n25570,
         n25571, n25572, n25573, n25574, n25575, n25576, n25577, n25578,
         n25579, n25580, n25581, n25582, n25583, n25584, n25585, n25586,
         n25587, n25588, n25589, n25590, n25591, n25592, n25593, n25594,
         n25595, n25596, n25597, n25598, n25599, n25600, n25601, n25602,
         n25603, n25604, n25605, n25606, n25607, n25608, n25609, n25610,
         n25611, n25612, n25613, n25614, n25615, n25616, n25617, n25618,
         n25619, n25620, n25621, n25622, n25623, n25624, n25625, n25626,
         n25627, n25628, n25629, n25630, n25631, n25632, n25633, n25634,
         n25635, n25636, n25637, n25638, n25639, n25640, n25641, n25642,
         n25643, n25644, n25645, n25646, n25647, n25648, n25649, n25650,
         n25651, n25652, n25653, n25654, n25655, n25656, n25657, n25658,
         n25659, n25660, n25661, n25662, n25663, n25664, n25665, n25666,
         n25667, n25668, n25669, n25670, n25671, n25672, n25673, n25674,
         n25675, n25676, n25677, n25678, n25679, n25680, n25681, n25682,
         n25683, n25684, n25685, n25686, n25687, n25688, n25689, n25690,
         n25691, n25692, n25693, n25694, n25695, n25696, n25697, n25698,
         n25699, n25700, n25701, n25702, n25703, n25704, n25705, n25706,
         n25707, n25708, n25709, n25710, n25711, n25712, n25713, n25714,
         n25715, n25716, n25717, n25718, n25719, n25720, n25721, n25722,
         n25723, n25724, n25725, n25726, n25727, n25728, n25729, n25730,
         n25731, n25732, n25733, n25734, n25735, n25736, n25737, n25738,
         n25739, n25740, n25741, n25742, n25743, n25744, n25745, n25746,
         n25747, n25748, n25749, n25750, n25751, n25752, n25753, n25754,
         n25755, n25756, n25757, n25758, n25759, n25760, n25761, n25762,
         n25763, n25764, n25765, n25766, n25767, n25768, n25769, n25770,
         n25771, n25772, n25773, n25774, n25775, n25776, n25777, n25778,
         n25779, n25780, n25781, n25782, n25783, n25784, n25785, n25786,
         n25787, n25788, n25789, n25790, n25791, n25792, n25793, n25794,
         n25795, n25796, n25797, n25798, n25799, n25800, n25801, n25802,
         n25803, n25804, n25805, n25806, n25807, n25808, n25809, n25810,
         n25811, n25812, n25813, n25814, n25815, n25816, n25817, n25818,
         n25819, n25820, n25821, n25822, n25823, n25824, n25825, n25826,
         n25827, n25828, n25829, n25830, n25831, n25832, n25833, n25834,
         n25835, n25836, n25837, n25838, n25839, n25840, n25841, n25842,
         n25843, n25844, n25845, n25846, n25847, n25848, n25849, n25850,
         n25851, n25852, n25853, n25854, n25855, n25856, n25857, n25858,
         n25859, n25860, n25861, n25862, n25863, n25864, n25865, n25866,
         n25867, n25868, n25869, n25870, n25871, n25872, n25873, n25874,
         n25875, n25876, n25877, n25878, n25879, n25880, n25881, n25882,
         n25883, n25884, n25885, n25886, n25887, n25888, n25889, n25890,
         n25891, n25892, n25893, n25894, n25895, n25896, n25897, n25898,
         n25899, n25900, n25901, n25902, n25903, n25904, n25905, n25906,
         n25907, n25908, n25909, n25910, n25911, n25912, n25913, n25914,
         n25915, n25916, n25917, n25918, n25919, n25920, n25921, n25922,
         n25923, n25924, n25925, n25926, n25927, n25928, n25929, n25930,
         n25931, n25932, n25933, n25934, n25935, n25936, n25937, n25938,
         n25939, n25940, n25941, n25942, n25943, n25944, n25945, n25946,
         n25947, n25948, n25949, n25950, n25951, n25952, n25953, n25954,
         n25955, n25956, n25957, n25958, n25959, n25960, n25961, n25962,
         n25963, n25964, n25965, n25966, n25967, n25968, n25969, n25970,
         n25971, n25972, n25973, n25974, n25975, n25976, n25977, n25978,
         n25979, n25980, n25981, n25982, n25983, n25984, n25985, n25986,
         n25987, n25988, n25989, n25990, n25991, n25992, n25993, n25994,
         n25995, n25996, n25997, n25998, n25999, n26000, n26001, n26002,
         n26003, n26004, n26005, n26006, n26007, n26008, n26009, n26010,
         n26011, n26012, n26013, n26014, n26015, n26016, n26017, n26018,
         n26019, n26020, n26021, n26022, n26023, n26024, n26025, n26026,
         n26027, n26028, n26029, n26030, n26031, n26032, n26033, n26034,
         n26035, n26036, n26037, n26038, n26039, n26040, n26041, n26042,
         n26043, n26044, n26045, n26046, n26047, n26048, n26049, n26050,
         n26051, n26052, n26053, n26054, n26055, n26056, n26057, n26058,
         n26059, n26060, n26061, n26062, n26063, n26064, n26065, n26066,
         n26067, n26068, n26069, n26070, n26071, n26072, n26073, n26074,
         n26075, n26076, n26077, n26078, n26079, n26080, n26081, n26082,
         n26083, n26084, n26085, n26086, n26087, n26088, n26089, n26090,
         n26091, n26092, n26093, n26094, n26095, n26096, n26097, n26098,
         n26099, n26100, n26101, n26102, n26103, n26104, n26105, n26106,
         n26107, n26108, n26109, n26110, n26111, n26112, n26113, n26114,
         n26115, n26116, n26117, n26118, n26119, n26120, n26121, n26122,
         n26123, n26124, n26125, n26126, n26127, n26128, n26129, n26130,
         n26131, n26132, n26133, n26134, n26135, n26136, n26137, n26138,
         n26139, n26140, n26141, n26142, n26143, n26144, n26145, n26146,
         n26147, n26148, n26149, n26150, n26151, n26152, n26153, n26154,
         n26155, n26156, n26157, n26158, n26159, n26160, n26161, n26162,
         n26163, n26164, n26165, n26166, n26167, n26168, n26169, n26170,
         n26171, n26172, n26173, n26174, n26175, n26176, n26177, n26178,
         n26179, n26180, n26181, n26182, n26183, n26184, n26185, n26186,
         n26187, n26188, n26189, n26190, n26191, n26192, n26193, n26194,
         n26195, n26196, n26197, n26198, n26199, n26200, n26201, n26202,
         n26203, n26204, n26205, n26206, n26207, n26208, n26209, n26210,
         n26211, n26212, n26213, n26214, n26215, n26216, n26217, n26218,
         n26219, n26220, n26221, n26222, n26223, n26224, n26225, n26226,
         n26227, n26228, n26229, n26230, n26231, n26232, n26233, n26234,
         n26235, n26236, n26237, n26238, n26239, n26240, n26241, n26242,
         n26243, n26244, n26245, n26246, n26247, n26248, n26249, n26250,
         n26251, n26252, n26253, n26254, n26255, n26256, n26257, n26258,
         n26259, n26260, n26261, n26262, n26263, n26264, n26265, n26266,
         n26267, n26268, n26269, n26270, n26271, n26272, n26273, n26274,
         n26275, n26276, n26277, n26278, n26279, n26280, n26281, n26282,
         n26283, n26284, n26285, n26286, n26287, n26288, n26289, n26290,
         n26291, n26292, n26293, n26294, n26295, n26296, n26297, n26298,
         n26299, n26300, n26301, n26302, n26303, n26304, n26305, n26306,
         n26307, n26308, n26309, n26310, n26311, n26312, n26313, n26314,
         n26315, n26316, n26317, n26318, n26319, n26320, n26321, n26322,
         n26323, n26324, n26325, n26326, n26327, n26328, n26329, n26330,
         n26331, n26332, n26333, n26334, n26335, n26336, n26337, n26338,
         n26339, n26340, n26341, n26342, n26343, n26344, n26345, n26346,
         n26347, n26348, n26349, n26350, n26351, n26352, n26353, n26354,
         n26355, n26356, n26357, n26358, n26359, n26360, n26361, n26362,
         n26363, n26364, n26365, n26366, n26367, n26368, n26369, n26370,
         n26371, n26372, n26373, n26374, n26375, n26376, n26377, n26378,
         n26379, n26380, n26381, n26382, n26383, n26384, n26385, n26386,
         n26387, n26388, n26389, n26390, n26391, n26392, n26393, n26394,
         n26395, n26396, n26397, n26398, n26399, n26400, n26401, n26402,
         n26403, n26404, n26405, n26406, n26407, n26408, n26409, n26410,
         n26411, n26412, n26413, n26414, n26415, n26416, n26417, n26418,
         n26419, n26420, n26421, n26422, n26423, n26424, n26425, n26426,
         n26427, n26428, n26429, n26430, n26431, n26432, n26433, n26434,
         n26435, n26436, n26437, n26438, n26439, n26440, n26441, n26442,
         n26443, n26444, n26445, n26446, n26447, n26448, n26449, n26450,
         n26451, n26452, n26453, n26454, n26455, n26456, n26457, n26458,
         n26459, n26460, n26461, n26462, n26463, n26464, n26465, n26466,
         n26467, n26468, n26469, n26470, n26471, n26472, n26473, n26474,
         n26475, n26476, n26477, n26478, n26479, n26480, n26481, n26482,
         n26483, n26484, n26485, n26486, n26487, n26488, n26489, n26490,
         n26491, n26492, n26493, n26494, n26495, n26496, n26497, n26498,
         n26499, n26500, n26501, n26502, n26503, n26504, n26505, n26506,
         n26507, n26508, n26509, n26510, n26511, n26512, n26513, n26514,
         n26515, n26516, n26517, n26518, n26519, n26520, n26521, n26522,
         n26523, n26524, n26525, n26526, n26527, n26528, n26529, n26530,
         n26531, n26532, n26533, n26534, n26535, n26536, n26537, n26538,
         n26539, n26540, n26541, n26542, n26543, n26544, n26545, n26546,
         n26547, n26548, n26549, n26550, n26551, n26552, n26553, n26554,
         n26555, n26556, n26557, n26558, n26559, n26560, n26561, n26562,
         n26563, n26564, n26565, n26566, n26567, n26568, n26569, n26570,
         n26571, n26572, n26573, n26574, n26575, n26576, n26577, n26578,
         n26579, n26580, n26581, n26582, n26583, n26584, n26585, n26586,
         n26587, n26588, n26589, n26590, n26591, n26592, n26593, n26594,
         n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602,
         n26603, n26604, n26605, n26606, n26607, n26608, n26609, n26610,
         n26611, n26612, n26613, n26614, n26615, n26616, n26617, n26618,
         n26619, n26620, n26621, n26622, n26623, n26624, n26625, n26626,
         n26627, n26628, n26629, n26630, n26631, n26632, n26633, n26634,
         n26635, n26636, n26637, n26638, n26639, n26640, n26641, n26642,
         n26643, n26644, n26645, n26646, n26647, n26648, n26649, n26650,
         n26651, n26652, n26653, n26654, n26655, n26656, n26657, n26658,
         n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666,
         n26667, n26668, n26669, n26670, n26671, n26672, n26673, n26674,
         n26675, n26676, n26677, n26678, n26679, n26680, n26681, n26682,
         n26683, n26684, n26685, n26686, n26687, n26688, n26689, n26690,
         n26691, n26692, n26693, n26694, n26695, n26696, n26697, n26698,
         n26699, n26700, n26701, n26702, n26703, n26704, n26705, n26706,
         n26707, n26708, n26709, n26710, n26711, n26712, n26713, n26714,
         n26715, n26716, n26717, n26718, n26719, n26720, n26721, n26722,
         n26723, n26724, n26725, n26726, n26727, n26728, n26729, n26730,
         n26731, n26732, n26733, n26734, n26735, n26736, n26737, n26738,
         n26739, n26740, n26741, n26742, n26743, n26744, n26745, n26746,
         n26747, n26748, n26749, n26750, n26751, n26752, n26753, n26754,
         n26755, n26756, n26757, n26758, n26759, n26760, n26761, n26762,
         n26763, n26764, n26765, n26766, n26767, n26768, n26769, n26770,
         n26771, n26772, n26773, n26774, n26775, n26776, n26777, n26778,
         n26779, n26780, n26781, n26782, n26783, n26784, n26785, n26786,
         n26787, n26788, n26789, n26790, n26791, n26792, n26793, n26794,
         n26795, n26796, n26797, n26798, n26799, n26800, n26801, n26802,
         n26803, n26804, n26805, n26806, n26807, n26808, n26809, n26810,
         n26811, n26812, n26813, n26814, n26815, n26816, n26817, n26818,
         n26819, n26820, n26821, n26822, n26823, n26824, n26825, n26826,
         n26827, n26828, n26829, n26830, n26831, n26832, n26833, n26834,
         n26835, n26836, n26837, n26838, n26839, n26840, n26841, n26842,
         n26843, n26844, n26845, n26846, n26847, n26848, n26849, n26850,
         n26851, n26852, n26853, n26854, n26855, n26856, n26857, n26858,
         n26859, n26860, n26861, n26862, n26863, n26864, n26865, n26866,
         n26867, n26868, n26869, n26870, n26871, n26872, n26873, n26874,
         n26875, n26876, n26877, n26878, n26879, n26880, n26881, n26882,
         n26883, n26884, n26885, n26886, n26887, n26888, n26889, n26890,
         n26891, n26892, n26893, n26894, n26895, n26896, n26897, n26898,
         n26899, n26900, n26901, n26902, n26903, n26904, n26905, n26906,
         n26907, n26908, n26909, n26910, n26911, n26912, n26913, n26914,
         n26915, n26916, n26917, n26918, n26919, n26920, n26921, n26922,
         n26923, n26924, n26925, n26926, n26927, n26928, n26929, n26930,
         n26931, n26932, n26933, n26934, n26935, n26936, n26937, n26938,
         n26939, n26940, n26941, n26942, n26943, n26944, n26945, n26946,
         n26947, n26948, n26949, n26950, n26951, n26952, n26953, n26954,
         n26955, n26956, n26957, n26958, n26959, n26960, n26961, n26962,
         n26963, n26964, n26965, n26966, n26967, n26968, n26969, n26970,
         n26971, n26972, n26973, n26974, n26975, n26976, n26977, n26978,
         n26979, n26980, n26981, n26982, n26983, n26984, n26985, n26986,
         n26987, n26988, n26989, n26990, n26991, n26992, n26993, n26994,
         n26995, n26996, n26997, n26998, n26999, n27000, n27001, n27002,
         n27003, n27004, n27005, n27006, n27007, n27008, n27009, n27010,
         n27011, n27012, n27013, n27014, n27015, n27016, n27017, n27018,
         n27019, n27020, n27021, n27022, n27023, n27024, n27025, n27026,
         n27027, n27028, n27029, n27030, n27031, n27032, n27033, n27034,
         n27035, n27036, n27037, n27038, n27039, n27040, n27041, n27042,
         n27043, n27044, n27045, n27046, n27047, n27048, n27049, n27050,
         n27051, n27052, n27053, n27054, n27055, n27056, n27057, n27058,
         n27059, n27060, n27061, n27062, n27063, n27064, n27065, n27066,
         n27067, n27068, n27069, n27070, n27071, n27072, n27073, n27074,
         n27075, n27076, n27077, n27078, n27079, n27080, n27081, n27082,
         n27083, n27084, n27085, n27086, n27087, n27088, n27089, n27090,
         n27091, n27092, n27093, n27094, n27095, n27096, n27097, n27098,
         n27099, n27100, n27101, n27102, n27103, n27104, n27105, n27106,
         n27107, n27108, n27109, n27110, n27111, n27112, n27113, n27114,
         n27115, n27116, n27117, n27118, n27119, n27120, n27121, n27122,
         n27123, n27124, n27125, n27126, n27127, n27128, n27129, n27130,
         n27131, n27132, n27133, n27134, n27135, n27136, n27137, n27138,
         n27139, n27140, n27141, n27142, n27143, n27144, n27145, n27146,
         n27147, n27148, n27149, n27150, n27151, n27152, n27153, n27154,
         n27155, n27156, n27157, n27158, n27159, n27160, n27161, n27162,
         n27163, n27164, n27165, n27166, n27167, n27168, n27169, n27170,
         n27171, n27172, n27173, n27174, n27175, n27176, n27177, n27178,
         n27179, n27180, n27181, n27182, n27183, n27184, n27185, n27186,
         n27187, n27188, n27189, n27190, n27191, n27192, n27193, n27194,
         n27195, n27196, n27197, n27198, n27199, n27200, n27201, n27202,
         n27203, n27204, n27205, n27206, n27207, n27208, n27209, n27210,
         n27211, n27212, n27213, n27214, n27215, n27216, n27217, n27218,
         n27219, n27220, n27221, n27222, n27223, n27224, n27225, n27226,
         n27227, n27228, n27229, n27230, n27231, n27232, n27233, n27234,
         n27235, n27236, n27237, n27238, n27239, n27240, n27241, n27242,
         n27243, n27244, n27245, n27246, n27247, n27248, n27249, n27250,
         n27251, n27252, n27253, n27254, n27255, n27256, n27257, n27258,
         n27259, n27260, n27261, n27262, n27263, n27264, n27265, n27266,
         n27267, n27268, n27269, n27270, n27271, n27272, n27273, n27274,
         n27275, n27276, n27277, n27278, n27279, n27280, n27281, n27282,
         n27283, n27284, n27285, n27286, n27287, n27288, n27289, n27290,
         n27291, n27292, n27293, n27294, n27295, n27296, n27297, n27298,
         n27299, n27300, n27301, n27302, n27303, n27304, n27305, n27306,
         n27307, n27308, n27309, n27310, n27311, n27312, n27313, n27314,
         n27315, n27316, n27317, n27318, n27319, n27320, n27321, n27322,
         n27323, n27324, n27325, n27326, n27327, n27328, n27329, n27330,
         n27331, n27332, n27333, n27334, n27335, n27336, n27337, n27338,
         n27339, n27340, n27341, n27342, n27343, n27344, n27345, n27346,
         n27347, n27348, n27349, n27350, n27351, n27352, n27353, n27354,
         n27355, n27356, n27357, n27358, n27359, n27360, n27361, n27362,
         n27363, n27364, n27365, n27366, n27367, n27368, n27369, n27370,
         n27371, n27372, n27373, n27374, n27375, n27376, n27377, n27378,
         n27379, n27380, n27381, n27382, n27383, n27384, n27385, n27386,
         n27387, n27388, n27389, n27390, n27391, n27392, n27393, n27394,
         n27395, n27396, n27397, n27398, n27399, n27400, n27401, n27402,
         n27403, n27404, n27405, n27406, n27407, n27408, n27409, n27410,
         n27411, n27412, n27413, n27414, n27415, n27416, n27417, n27418,
         n27419, n27420, n27421, n27422, n27423, n27424, n27425, n27426,
         n27427, n27428, n27429, n27430, n27431, n27432, n27433, n27434,
         n27435, n27436, n27437, n27438, n27439, n27440, n27441, n27442,
         n27443, n27444, n27445, n27446, n27447, n27448, n27449, n27450,
         n27451, n27452, n27453, n27454, n27455, n27456, n27457, n27458,
         n27459, n27460, n27461, n27462, n27463, n27464, n27465, n27466,
         n27467, n27468, n27469, n27470, n27471, n27472, n27473, n27474,
         n27475, n27476, n27477, n27478, n27479, n27480, n27481, n27482,
         n27483, n27484, n27485, n27486, n27487, n27488, n27489, n27490,
         n27491, n27492, n27493, n27494, n27495, n27496, n27497, n27498,
         n27499, n27500, n27501, n27502, n27503, n27504, n27505, n27506,
         n27507, n27508, n27509, n27510, n27511, n27512, n27513, n27514,
         n27515, n27516, n27517, n27518, n27519, n27520, n27521, n27522,
         n27523, n27524, n27525, n27526, n27527, n27528, n27529, n27530,
         n27531, n27532, n27533, n27534, n27535, n27536, n27537, n27538,
         n27539, n27540, n27541, n27542, n27543, n27544, n27545, n27546,
         n27547, n27548, n27549, n27550, n27551, n27552, n27553, n27554,
         n27555, n27556, n27557, n27558, n27559, n27560, n27561, n27562,
         n27563, n27564, n27565, n27566, n27567, n27568, n27569, n27570,
         n27571, n27572, n27573, n27574, n27575, n27576, n27577, n27578,
         n27579, n27580, n27581, n27582, n27583, n27584, n27585, n27586,
         n27587, n27588, n27589, n27590, n27591, n27592;

  dp_1 \x_reg[120][15]  ( .ip(n17322), .ck(clk), .q(\x[120][15] ) );
  dp_1 \x_reg[120][14]  ( .ip(n17321), .ck(clk), .q(\x[120][14] ) );
  dp_1 \x_reg[120][13]  ( .ip(n17320), .ck(clk), .q(\x[120][13] ) );
  dp_1 \x_reg[120][12]  ( .ip(n17319), .ck(clk), .q(\x[120][12] ) );
  dp_1 \x_reg[120][11]  ( .ip(n17318), .ck(clk), .q(\x[120][11] ) );
  dp_1 \x_reg[120][10]  ( .ip(n17317), .ck(clk), .q(\x[120][10] ) );
  dp_1 \x_reg[120][9]  ( .ip(n17316), .ck(clk), .q(\x[120][9] ) );
  dp_1 \x_reg[120][8]  ( .ip(n17315), .ck(clk), .q(\x[120][8] ) );
  dp_1 \x_reg[120][7]  ( .ip(n17314), .ck(clk), .q(\x[120][7] ) );
  dp_1 \x_reg[120][6]  ( .ip(n17313), .ck(clk), .q(\x[120][6] ) );
  dp_1 \x_reg[120][5]  ( .ip(n17312), .ck(clk), .q(\x[120][5] ) );
  dp_1 \x_reg[120][4]  ( .ip(n17311), .ck(clk), .q(\x[120][4] ) );
  dp_1 \x_reg[120][3]  ( .ip(n17310), .ck(clk), .q(\x[120][3] ) );
  dp_1 \x_reg[120][2]  ( .ip(n17309), .ck(clk), .q(\x[120][2] ) );
  dp_1 \x_reg[120][1]  ( .ip(n17308), .ck(clk), .q(\x[120][1] ) );
  dp_1 \x_reg[120][0]  ( .ip(n17307), .ck(clk), .q(\x[120][0] ) );
  dp_1 \x_reg[119][15]  ( .ip(n17306), .ck(clk), .q(\x[119][15] ) );
  dp_1 \x_reg[119][14]  ( .ip(n17305), .ck(clk), .q(\x[119][14] ) );
  dp_1 \x_reg[119][13]  ( .ip(n17304), .ck(clk), .q(\x[119][13] ) );
  dp_1 \x_reg[119][12]  ( .ip(n17303), .ck(clk), .q(\x[119][12] ) );
  dp_1 \x_reg[119][11]  ( .ip(n17302), .ck(clk), .q(\x[119][11] ) );
  dp_1 \x_reg[119][10]  ( .ip(n17301), .ck(clk), .q(\x[119][10] ) );
  dp_1 \x_reg[119][9]  ( .ip(n17300), .ck(clk), .q(\x[119][9] ) );
  dp_1 \x_reg[119][8]  ( .ip(n17299), .ck(clk), .q(\x[119][8] ) );
  dp_1 \x_reg[119][7]  ( .ip(n17298), .ck(clk), .q(\x[119][7] ) );
  dp_1 \x_reg[119][6]  ( .ip(n17297), .ck(clk), .q(\x[119][6] ) );
  dp_1 \x_reg[119][5]  ( .ip(n17296), .ck(clk), .q(\x[119][5] ) );
  dp_1 \x_reg[119][4]  ( .ip(n17295), .ck(clk), .q(\x[119][4] ) );
  dp_1 \x_reg[119][3]  ( .ip(n17294), .ck(clk), .q(\x[119][3] ) );
  dp_1 \x_reg[119][2]  ( .ip(n17293), .ck(clk), .q(\x[119][2] ) );
  dp_1 \x_reg[119][1]  ( .ip(n17292), .ck(clk), .q(\x[119][1] ) );
  dp_1 \x_reg[119][0]  ( .ip(n17291), .ck(clk), .q(\x[119][0] ) );
  dp_1 \x_reg[118][15]  ( .ip(n17290), .ck(clk), .q(\x[118][15] ) );
  dp_1 \x_reg[118][14]  ( .ip(n17289), .ck(clk), .q(\x[118][14] ) );
  dp_1 \x_reg[118][13]  ( .ip(n17288), .ck(clk), .q(\x[118][13] ) );
  dp_1 \x_reg[118][12]  ( .ip(n17287), .ck(clk), .q(\x[118][12] ) );
  dp_1 \x_reg[118][11]  ( .ip(n17286), .ck(clk), .q(\x[118][11] ) );
  dp_1 \x_reg[118][10]  ( .ip(n17285), .ck(clk), .q(\x[118][10] ) );
  dp_1 \x_reg[118][9]  ( .ip(n17284), .ck(clk), .q(\x[118][9] ) );
  dp_1 \x_reg[118][8]  ( .ip(n17283), .ck(clk), .q(\x[118][8] ) );
  dp_1 \x_reg[118][7]  ( .ip(n17282), .ck(clk), .q(\x[118][7] ) );
  dp_1 \x_reg[118][6]  ( .ip(n17281), .ck(clk), .q(\x[118][6] ) );
  dp_1 \x_reg[118][5]  ( .ip(n17280), .ck(clk), .q(\x[118][5] ) );
  dp_1 \x_reg[118][4]  ( .ip(n17279), .ck(clk), .q(\x[118][4] ) );
  dp_1 \x_reg[118][3]  ( .ip(n17278), .ck(clk), .q(\x[118][3] ) );
  dp_1 \x_reg[118][2]  ( .ip(n17277), .ck(clk), .q(\x[118][2] ) );
  dp_1 \x_reg[118][1]  ( .ip(n17276), .ck(clk), .q(\x[118][1] ) );
  dp_1 \x_reg[118][0]  ( .ip(n17275), .ck(clk), .q(\x[118][0] ) );
  dp_1 \x_reg[117][15]  ( .ip(n17274), .ck(clk), .q(\x[117][15] ) );
  dp_1 \x_reg[117][14]  ( .ip(n17273), .ck(clk), .q(\x[117][14] ) );
  dp_1 \x_reg[117][13]  ( .ip(n17272), .ck(clk), .q(\x[117][13] ) );
  dp_1 \x_reg[117][12]  ( .ip(n17271), .ck(clk), .q(\x[117][12] ) );
  dp_1 \x_reg[117][11]  ( .ip(n17270), .ck(clk), .q(\x[117][11] ) );
  dp_1 \x_reg[117][10]  ( .ip(n17269), .ck(clk), .q(\x[117][10] ) );
  dp_1 \x_reg[117][9]  ( .ip(n17268), .ck(clk), .q(\x[117][9] ) );
  dp_1 \x_reg[117][8]  ( .ip(n17267), .ck(clk), .q(\x[117][8] ) );
  dp_1 \x_reg[117][7]  ( .ip(n17266), .ck(clk), .q(\x[117][7] ) );
  dp_1 \x_reg[117][6]  ( .ip(n17265), .ck(clk), .q(\x[117][6] ) );
  dp_1 \x_reg[117][5]  ( .ip(n17264), .ck(clk), .q(\x[117][5] ) );
  dp_1 \x_reg[117][4]  ( .ip(n17263), .ck(clk), .q(\x[117][4] ) );
  dp_1 \x_reg[117][3]  ( .ip(n17262), .ck(clk), .q(\x[117][3] ) );
  dp_1 \x_reg[117][2]  ( .ip(n17261), .ck(clk), .q(\x[117][2] ) );
  dp_1 \x_reg[117][1]  ( .ip(n17260), .ck(clk), .q(\x[117][1] ) );
  dp_1 \x_reg[117][0]  ( .ip(n17259), .ck(clk), .q(\x[117][0] ) );
  dp_1 \x_reg[116][15]  ( .ip(n17258), .ck(clk), .q(\x[116][15] ) );
  dp_1 \x_reg[116][14]  ( .ip(n17257), .ck(clk), .q(\x[116][14] ) );
  dp_1 \x_reg[116][13]  ( .ip(n17256), .ck(clk), .q(\x[116][13] ) );
  dp_1 \x_reg[116][12]  ( .ip(n17255), .ck(clk), .q(\x[116][12] ) );
  dp_1 \x_reg[116][11]  ( .ip(n17254), .ck(clk), .q(\x[116][11] ) );
  dp_1 \x_reg[116][10]  ( .ip(n17253), .ck(clk), .q(\x[116][10] ) );
  dp_1 \x_reg[116][9]  ( .ip(n17252), .ck(clk), .q(\x[116][9] ) );
  dp_1 \x_reg[116][8]  ( .ip(n17251), .ck(clk), .q(\x[116][8] ) );
  dp_1 \x_reg[116][7]  ( .ip(n17250), .ck(clk), .q(\x[116][7] ) );
  dp_1 \x_reg[116][6]  ( .ip(n17249), .ck(clk), .q(\x[116][6] ) );
  dp_1 \x_reg[116][5]  ( .ip(n17248), .ck(clk), .q(\x[116][5] ) );
  dp_1 \x_reg[116][4]  ( .ip(n17247), .ck(clk), .q(\x[116][4] ) );
  dp_1 \x_reg[116][3]  ( .ip(n17246), .ck(clk), .q(\x[116][3] ) );
  dp_1 \x_reg[116][2]  ( .ip(n17245), .ck(clk), .q(\x[116][2] ) );
  dp_1 \x_reg[116][1]  ( .ip(n17244), .ck(clk), .q(\x[116][1] ) );
  dp_1 \x_reg[116][0]  ( .ip(n17243), .ck(clk), .q(\x[116][0] ) );
  dp_1 \x_reg[115][15]  ( .ip(n17242), .ck(clk), .q(\x[115][15] ) );
  dp_1 \x_reg[115][14]  ( .ip(n17241), .ck(clk), .q(\x[115][14] ) );
  dp_1 \x_reg[115][13]  ( .ip(n17240), .ck(clk), .q(\x[115][13] ) );
  dp_1 \x_reg[115][12]  ( .ip(n17239), .ck(clk), .q(\x[115][12] ) );
  dp_1 \x_reg[115][11]  ( .ip(n17238), .ck(clk), .q(\x[115][11] ) );
  dp_1 \x_reg[115][10]  ( .ip(n17237), .ck(clk), .q(\x[115][10] ) );
  dp_1 \x_reg[115][9]  ( .ip(n17236), .ck(clk), .q(\x[115][9] ) );
  dp_1 \x_reg[115][8]  ( .ip(n17235), .ck(clk), .q(\x[115][8] ) );
  dp_1 \x_reg[115][7]  ( .ip(n17234), .ck(clk), .q(\x[115][7] ) );
  dp_1 \x_reg[115][6]  ( .ip(n17233), .ck(clk), .q(\x[115][6] ) );
  dp_1 \x_reg[115][5]  ( .ip(n17232), .ck(clk), .q(\x[115][5] ) );
  dp_1 \x_reg[115][4]  ( .ip(n17231), .ck(clk), .q(\x[115][4] ) );
  dp_1 \x_reg[115][3]  ( .ip(n17230), .ck(clk), .q(\x[115][3] ) );
  dp_1 \x_reg[115][2]  ( .ip(n17229), .ck(clk), .q(\x[115][2] ) );
  dp_1 \x_reg[115][1]  ( .ip(n17228), .ck(clk), .q(\x[115][1] ) );
  dp_1 \x_reg[115][0]  ( .ip(n17227), .ck(clk), .q(\x[115][0] ) );
  dp_1 \x_reg[114][15]  ( .ip(n17226), .ck(clk), .q(\x[114][15] ) );
  dp_1 \x_reg[114][14]  ( .ip(n17225), .ck(clk), .q(\x[114][14] ) );
  dp_1 \x_reg[114][13]  ( .ip(n17224), .ck(clk), .q(\x[114][13] ) );
  dp_1 \x_reg[114][12]  ( .ip(n17223), .ck(clk), .q(\x[114][12] ) );
  dp_1 \x_reg[114][11]  ( .ip(n17222), .ck(clk), .q(\x[114][11] ) );
  dp_1 \x_reg[114][10]  ( .ip(n17221), .ck(clk), .q(\x[114][10] ) );
  dp_1 \x_reg[114][9]  ( .ip(n17220), .ck(clk), .q(\x[114][9] ) );
  dp_1 \x_reg[114][8]  ( .ip(n17219), .ck(clk), .q(\x[114][8] ) );
  dp_1 \x_reg[114][7]  ( .ip(n17218), .ck(clk), .q(\x[114][7] ) );
  dp_1 \x_reg[114][6]  ( .ip(n17217), .ck(clk), .q(\x[114][6] ) );
  dp_1 \x_reg[114][5]  ( .ip(n17216), .ck(clk), .q(\x[114][5] ) );
  dp_1 \x_reg[114][4]  ( .ip(n17215), .ck(clk), .q(\x[114][4] ) );
  dp_1 \x_reg[114][3]  ( .ip(n17214), .ck(clk), .q(\x[114][3] ) );
  dp_1 \x_reg[114][2]  ( .ip(n17213), .ck(clk), .q(\x[114][2] ) );
  dp_1 \x_reg[114][1]  ( .ip(n17212), .ck(clk), .q(\x[114][1] ) );
  dp_1 \x_reg[114][0]  ( .ip(n17211), .ck(clk), .q(\x[114][0] ) );
  dp_1 \x_reg[113][15]  ( .ip(n17210), .ck(clk), .q(\x[113][15] ) );
  dp_1 \x_reg[113][14]  ( .ip(n17209), .ck(clk), .q(\x[113][14] ) );
  dp_1 \x_reg[113][13]  ( .ip(n17208), .ck(clk), .q(\x[113][13] ) );
  dp_1 \x_reg[113][12]  ( .ip(n17207), .ck(clk), .q(\x[113][12] ) );
  dp_1 \x_reg[113][11]  ( .ip(n17206), .ck(clk), .q(\x[113][11] ) );
  dp_1 \x_reg[113][10]  ( .ip(n17205), .ck(clk), .q(\x[113][10] ) );
  dp_1 \x_reg[113][9]  ( .ip(n17204), .ck(clk), .q(\x[113][9] ) );
  dp_1 \x_reg[113][8]  ( .ip(n17203), .ck(clk), .q(\x[113][8] ) );
  dp_1 \x_reg[113][7]  ( .ip(n17202), .ck(clk), .q(\x[113][7] ) );
  dp_1 \x_reg[113][6]  ( .ip(n17201), .ck(clk), .q(\x[113][6] ) );
  dp_1 \x_reg[113][5]  ( .ip(n17200), .ck(clk), .q(\x[113][5] ) );
  dp_1 \x_reg[113][4]  ( .ip(n17199), .ck(clk), .q(\x[113][4] ) );
  dp_1 \x_reg[113][3]  ( .ip(n17198), .ck(clk), .q(\x[113][3] ) );
  dp_1 \x_reg[113][2]  ( .ip(n17197), .ck(clk), .q(\x[113][2] ) );
  dp_1 \x_reg[113][1]  ( .ip(n17196), .ck(clk), .q(\x[113][1] ) );
  dp_1 \x_reg[113][0]  ( .ip(n17195), .ck(clk), .q(\x[113][0] ) );
  dp_1 \x_reg[112][15]  ( .ip(n17194), .ck(clk), .q(\x[112][15] ) );
  dp_1 \x_reg[112][14]  ( .ip(n17193), .ck(clk), .q(\x[112][14] ) );
  dp_1 \x_reg[112][13]  ( .ip(n17192), .ck(clk), .q(\x[112][13] ) );
  dp_1 \x_reg[112][12]  ( .ip(n17191), .ck(clk), .q(\x[112][12] ) );
  dp_1 \x_reg[112][11]  ( .ip(n17190), .ck(clk), .q(\x[112][11] ) );
  dp_1 \x_reg[112][10]  ( .ip(n17189), .ck(clk), .q(\x[112][10] ) );
  dp_1 \x_reg[112][9]  ( .ip(n17188), .ck(clk), .q(\x[112][9] ) );
  dp_1 \x_reg[112][8]  ( .ip(n17187), .ck(clk), .q(\x[112][8] ) );
  dp_1 \x_reg[112][7]  ( .ip(n17186), .ck(clk), .q(\x[112][7] ) );
  dp_1 \x_reg[112][6]  ( .ip(n17185), .ck(clk), .q(\x[112][6] ) );
  dp_1 \x_reg[112][5]  ( .ip(n17184), .ck(clk), .q(\x[112][5] ) );
  dp_1 \x_reg[112][4]  ( .ip(n17183), .ck(clk), .q(\x[112][4] ) );
  dp_1 \x_reg[112][3]  ( .ip(n17182), .ck(clk), .q(\x[112][3] ) );
  dp_1 \x_reg[112][2]  ( .ip(n17181), .ck(clk), .q(\x[112][2] ) );
  dp_1 \x_reg[112][1]  ( .ip(n17180), .ck(clk), .q(\x[112][1] ) );
  dp_1 \x_reg[112][0]  ( .ip(n17179), .ck(clk), .q(\x[112][0] ) );
  dp_1 \x_reg[111][15]  ( .ip(n17178), .ck(clk), .q(\x[111][15] ) );
  dp_1 \x_reg[111][14]  ( .ip(n17177), .ck(clk), .q(\x[111][14] ) );
  dp_1 \x_reg[111][13]  ( .ip(n17176), .ck(clk), .q(\x[111][13] ) );
  dp_1 \x_reg[111][12]  ( .ip(n17175), .ck(clk), .q(\x[111][12] ) );
  dp_1 \x_reg[111][11]  ( .ip(n17174), .ck(clk), .q(\x[111][11] ) );
  dp_1 \x_reg[111][10]  ( .ip(n17173), .ck(clk), .q(\x[111][10] ) );
  dp_1 \x_reg[111][9]  ( .ip(n17172), .ck(clk), .q(\x[111][9] ) );
  dp_1 \x_reg[111][8]  ( .ip(n17171), .ck(clk), .q(\x[111][8] ) );
  dp_1 \x_reg[111][7]  ( .ip(n17170), .ck(clk), .q(\x[111][7] ) );
  dp_1 \x_reg[111][6]  ( .ip(n17169), .ck(clk), .q(\x[111][6] ) );
  dp_1 \x_reg[111][5]  ( .ip(n17168), .ck(clk), .q(\x[111][5] ) );
  dp_1 \x_reg[111][4]  ( .ip(n17167), .ck(clk), .q(\x[111][4] ) );
  dp_1 \x_reg[111][3]  ( .ip(n17166), .ck(clk), .q(\x[111][3] ) );
  dp_1 \x_reg[111][2]  ( .ip(n17165), .ck(clk), .q(\x[111][2] ) );
  dp_1 \x_reg[111][1]  ( .ip(n17164), .ck(clk), .q(\x[111][1] ) );
  dp_1 \x_reg[111][0]  ( .ip(n17163), .ck(clk), .q(\x[111][0] ) );
  dp_1 \x_reg[110][15]  ( .ip(n17162), .ck(clk), .q(\x[110][15] ) );
  dp_1 \x_reg[110][14]  ( .ip(n17161), .ck(clk), .q(\x[110][14] ) );
  dp_1 \x_reg[110][13]  ( .ip(n17160), .ck(clk), .q(\x[110][13] ) );
  dp_1 \x_reg[110][12]  ( .ip(n17159), .ck(clk), .q(\x[110][12] ) );
  dp_1 \x_reg[110][11]  ( .ip(n17158), .ck(clk), .q(\x[110][11] ) );
  dp_1 \x_reg[110][10]  ( .ip(n17157), .ck(clk), .q(\x[110][10] ) );
  dp_1 \x_reg[110][9]  ( .ip(n17156), .ck(clk), .q(\x[110][9] ) );
  dp_1 \x_reg[110][8]  ( .ip(n17155), .ck(clk), .q(\x[110][8] ) );
  dp_1 \x_reg[110][7]  ( .ip(n17154), .ck(clk), .q(\x[110][7] ) );
  dp_1 \x_reg[110][6]  ( .ip(n17153), .ck(clk), .q(\x[110][6] ) );
  dp_1 \x_reg[110][5]  ( .ip(n17152), .ck(clk), .q(\x[110][5] ) );
  dp_1 \x_reg[110][4]  ( .ip(n17151), .ck(clk), .q(\x[110][4] ) );
  dp_1 \x_reg[110][3]  ( .ip(n17150), .ck(clk), .q(\x[110][3] ) );
  dp_1 \x_reg[110][2]  ( .ip(n17149), .ck(clk), .q(\x[110][2] ) );
  dp_1 \x_reg[110][1]  ( .ip(n17148), .ck(clk), .q(\x[110][1] ) );
  dp_1 \x_reg[110][0]  ( .ip(n17147), .ck(clk), .q(\x[110][0] ) );
  dp_1 \x_reg[109][15]  ( .ip(n17146), .ck(clk), .q(\x[109][15] ) );
  dp_1 \x_reg[109][14]  ( .ip(n17145), .ck(clk), .q(\x[109][14] ) );
  dp_1 \x_reg[109][13]  ( .ip(n17144), .ck(clk), .q(\x[109][13] ) );
  dp_1 \x_reg[109][12]  ( .ip(n17143), .ck(clk), .q(\x[109][12] ) );
  dp_1 \x_reg[109][11]  ( .ip(n17142), .ck(clk), .q(\x[109][11] ) );
  dp_1 \x_reg[109][10]  ( .ip(n17141), .ck(clk), .q(\x[109][10] ) );
  dp_1 \x_reg[109][9]  ( .ip(n17140), .ck(clk), .q(\x[109][9] ) );
  dp_1 \x_reg[109][8]  ( .ip(n17139), .ck(clk), .q(\x[109][8] ) );
  dp_1 \x_reg[109][7]  ( .ip(n17138), .ck(clk), .q(\x[109][7] ) );
  dp_1 \x_reg[109][6]  ( .ip(n17137), .ck(clk), .q(\x[109][6] ) );
  dp_1 \x_reg[109][5]  ( .ip(n17136), .ck(clk), .q(\x[109][5] ) );
  dp_1 \x_reg[109][4]  ( .ip(n17135), .ck(clk), .q(\x[109][4] ) );
  dp_1 \x_reg[109][3]  ( .ip(n17134), .ck(clk), .q(\x[109][3] ) );
  dp_1 \x_reg[109][2]  ( .ip(n17133), .ck(clk), .q(\x[109][2] ) );
  dp_1 \x_reg[109][1]  ( .ip(n17132), .ck(clk), .q(\x[109][1] ) );
  dp_1 \x_reg[109][0]  ( .ip(n17131), .ck(clk), .q(\x[109][0] ) );
  dp_1 \x_reg[108][15]  ( .ip(n17130), .ck(clk), .q(\x[108][15] ) );
  dp_1 \x_reg[108][14]  ( .ip(n17129), .ck(clk), .q(\x[108][14] ) );
  dp_1 \x_reg[108][13]  ( .ip(n17128), .ck(clk), .q(\x[108][13] ) );
  dp_1 \x_reg[108][12]  ( .ip(n17127), .ck(clk), .q(\x[108][12] ) );
  dp_1 \x_reg[108][11]  ( .ip(n17126), .ck(clk), .q(\x[108][11] ) );
  dp_1 \x_reg[108][10]  ( .ip(n17125), .ck(clk), .q(\x[108][10] ) );
  dp_1 \x_reg[108][9]  ( .ip(n17124), .ck(clk), .q(\x[108][9] ) );
  dp_1 \x_reg[108][8]  ( .ip(n17123), .ck(clk), .q(\x[108][8] ) );
  dp_1 \x_reg[108][7]  ( .ip(n17122), .ck(clk), .q(\x[108][7] ) );
  dp_1 \x_reg[108][6]  ( .ip(n17121), .ck(clk), .q(\x[108][6] ) );
  dp_1 \x_reg[108][5]  ( .ip(n17120), .ck(clk), .q(\x[108][5] ) );
  dp_1 \x_reg[108][4]  ( .ip(n17119), .ck(clk), .q(\x[108][4] ) );
  dp_1 \x_reg[108][3]  ( .ip(n17118), .ck(clk), .q(\x[108][3] ) );
  dp_1 \x_reg[108][2]  ( .ip(n17117), .ck(clk), .q(\x[108][2] ) );
  dp_1 \x_reg[108][1]  ( .ip(n17116), .ck(clk), .q(\x[108][1] ) );
  dp_1 \x_reg[108][0]  ( .ip(n17115), .ck(clk), .q(\x[108][0] ) );
  dp_1 \x_reg[107][15]  ( .ip(n17114), .ck(clk), .q(\x[107][15] ) );
  dp_1 \x_reg[107][14]  ( .ip(n17113), .ck(clk), .q(\x[107][14] ) );
  dp_1 \x_reg[107][13]  ( .ip(n17112), .ck(clk), .q(\x[107][13] ) );
  dp_1 \x_reg[107][12]  ( .ip(n17111), .ck(clk), .q(\x[107][12] ) );
  dp_1 \x_reg[107][11]  ( .ip(n17110), .ck(clk), .q(\x[107][11] ) );
  dp_1 \x_reg[107][10]  ( .ip(n17109), .ck(clk), .q(\x[107][10] ) );
  dp_1 \x_reg[107][9]  ( .ip(n17108), .ck(clk), .q(\x[107][9] ) );
  dp_1 \x_reg[107][8]  ( .ip(n17107), .ck(clk), .q(\x[107][8] ) );
  dp_1 \x_reg[107][7]  ( .ip(n17106), .ck(clk), .q(\x[107][7] ) );
  dp_1 \x_reg[107][6]  ( .ip(n17105), .ck(clk), .q(\x[107][6] ) );
  dp_1 \x_reg[107][5]  ( .ip(n17104), .ck(clk), .q(\x[107][5] ) );
  dp_1 \x_reg[107][4]  ( .ip(n17103), .ck(clk), .q(\x[107][4] ) );
  dp_1 \x_reg[107][3]  ( .ip(n17102), .ck(clk), .q(\x[107][3] ) );
  dp_1 \x_reg[107][2]  ( .ip(n17101), .ck(clk), .q(\x[107][2] ) );
  dp_1 \x_reg[107][1]  ( .ip(n17100), .ck(clk), .q(\x[107][1] ) );
  dp_1 \x_reg[107][0]  ( .ip(n17099), .ck(clk), .q(\x[107][0] ) );
  dp_1 \x_reg[106][15]  ( .ip(n17098), .ck(clk), .q(\x[106][15] ) );
  dp_1 \x_reg[106][14]  ( .ip(n17097), .ck(clk), .q(\x[106][14] ) );
  dp_1 \x_reg[106][13]  ( .ip(n17096), .ck(clk), .q(\x[106][13] ) );
  dp_1 \x_reg[106][12]  ( .ip(n17095), .ck(clk), .q(\x[106][12] ) );
  dp_1 \x_reg[106][11]  ( .ip(n17094), .ck(clk), .q(\x[106][11] ) );
  dp_1 \x_reg[106][10]  ( .ip(n17093), .ck(clk), .q(\x[106][10] ) );
  dp_1 \x_reg[106][9]  ( .ip(n17092), .ck(clk), .q(\x[106][9] ) );
  dp_1 \x_reg[106][8]  ( .ip(n17091), .ck(clk), .q(\x[106][8] ) );
  dp_1 \x_reg[106][7]  ( .ip(n17090), .ck(clk), .q(\x[106][7] ) );
  dp_1 \x_reg[106][6]  ( .ip(n17089), .ck(clk), .q(\x[106][6] ) );
  dp_1 \x_reg[106][5]  ( .ip(n17088), .ck(clk), .q(\x[106][5] ) );
  dp_1 \x_reg[106][4]  ( .ip(n17087), .ck(clk), .q(\x[106][4] ) );
  dp_1 \x_reg[106][3]  ( .ip(n17086), .ck(clk), .q(\x[106][3] ) );
  dp_1 \x_reg[106][2]  ( .ip(n17085), .ck(clk), .q(\x[106][2] ) );
  dp_1 \x_reg[106][1]  ( .ip(n17084), .ck(clk), .q(\x[106][1] ) );
  dp_1 \x_reg[106][0]  ( .ip(n17083), .ck(clk), .q(\x[106][0] ) );
  dp_1 \x_reg[105][15]  ( .ip(n17082), .ck(clk), .q(\x[105][15] ) );
  dp_1 \x_reg[105][14]  ( .ip(n17081), .ck(clk), .q(\x[105][14] ) );
  dp_1 \x_reg[105][13]  ( .ip(n17080), .ck(clk), .q(\x[105][13] ) );
  dp_1 \x_reg[105][12]  ( .ip(n17079), .ck(clk), .q(\x[105][12] ) );
  dp_1 \x_reg[105][11]  ( .ip(n17078), .ck(clk), .q(\x[105][11] ) );
  dp_1 \x_reg[105][10]  ( .ip(n17077), .ck(clk), .q(\x[105][10] ) );
  dp_1 \x_reg[105][9]  ( .ip(n17076), .ck(clk), .q(\x[105][9] ) );
  dp_1 \x_reg[105][8]  ( .ip(n17075), .ck(clk), .q(\x[105][8] ) );
  dp_1 \x_reg[105][7]  ( .ip(n17074), .ck(clk), .q(\x[105][7] ) );
  dp_1 \x_reg[105][6]  ( .ip(n17073), .ck(clk), .q(\x[105][6] ) );
  dp_1 \x_reg[105][5]  ( .ip(n17072), .ck(clk), .q(\x[105][5] ) );
  dp_1 \x_reg[105][4]  ( .ip(n17071), .ck(clk), .q(\x[105][4] ) );
  dp_1 \x_reg[105][3]  ( .ip(n17070), .ck(clk), .q(\x[105][3] ) );
  dp_1 \x_reg[105][2]  ( .ip(n17069), .ck(clk), .q(\x[105][2] ) );
  dp_1 \x_reg[105][1]  ( .ip(n17068), .ck(clk), .q(\x[105][1] ) );
  dp_1 \x_reg[105][0]  ( .ip(n17067), .ck(clk), .q(\x[105][0] ) );
  dp_1 \x_reg[104][15]  ( .ip(n17066), .ck(clk), .q(\x[104][15] ) );
  dp_1 \x_reg[104][14]  ( .ip(n17065), .ck(clk), .q(\x[104][14] ) );
  dp_1 \x_reg[104][13]  ( .ip(n17064), .ck(clk), .q(\x[104][13] ) );
  dp_1 \x_reg[104][12]  ( .ip(n17063), .ck(clk), .q(\x[104][12] ) );
  dp_1 \x_reg[104][11]  ( .ip(n17062), .ck(clk), .q(\x[104][11] ) );
  dp_1 \x_reg[104][10]  ( .ip(n17061), .ck(clk), .q(\x[104][10] ) );
  dp_1 \x_reg[104][9]  ( .ip(n17060), .ck(clk), .q(\x[104][9] ) );
  dp_1 \x_reg[104][8]  ( .ip(n17059), .ck(clk), .q(\x[104][8] ) );
  dp_1 \x_reg[104][7]  ( .ip(n17058), .ck(clk), .q(\x[104][7] ) );
  dp_1 \x_reg[104][6]  ( .ip(n17057), .ck(clk), .q(\x[104][6] ) );
  dp_1 \x_reg[104][5]  ( .ip(n17056), .ck(clk), .q(\x[104][5] ) );
  dp_1 \x_reg[104][4]  ( .ip(n17055), .ck(clk), .q(\x[104][4] ) );
  dp_1 \x_reg[104][3]  ( .ip(n17054), .ck(clk), .q(\x[104][3] ) );
  dp_1 \x_reg[104][2]  ( .ip(n17053), .ck(clk), .q(\x[104][2] ) );
  dp_1 \x_reg[104][1]  ( .ip(n17052), .ck(clk), .q(\x[104][1] ) );
  dp_1 \x_reg[104][0]  ( .ip(n17051), .ck(clk), .q(\x[104][0] ) );
  dp_1 \x_reg[103][15]  ( .ip(n17050), .ck(clk), .q(\x[103][15] ) );
  dp_1 \x_reg[103][14]  ( .ip(n17049), .ck(clk), .q(\x[103][14] ) );
  dp_1 \x_reg[103][13]  ( .ip(n17048), .ck(clk), .q(\x[103][13] ) );
  dp_1 \x_reg[103][12]  ( .ip(n17047), .ck(clk), .q(\x[103][12] ) );
  dp_1 \x_reg[103][11]  ( .ip(n17046), .ck(clk), .q(\x[103][11] ) );
  dp_1 \x_reg[103][10]  ( .ip(n17045), .ck(clk), .q(\x[103][10] ) );
  dp_1 \x_reg[103][9]  ( .ip(n17044), .ck(clk), .q(\x[103][9] ) );
  dp_1 \x_reg[103][8]  ( .ip(n17043), .ck(clk), .q(\x[103][8] ) );
  dp_1 \x_reg[103][7]  ( .ip(n17042), .ck(clk), .q(\x[103][7] ) );
  dp_1 \x_reg[103][6]  ( .ip(n17041), .ck(clk), .q(\x[103][6] ) );
  dp_1 \x_reg[103][5]  ( .ip(n17040), .ck(clk), .q(\x[103][5] ) );
  dp_1 \x_reg[103][4]  ( .ip(n17039), .ck(clk), .q(\x[103][4] ) );
  dp_1 \x_reg[103][3]  ( .ip(n17038), .ck(clk), .q(\x[103][3] ) );
  dp_1 \x_reg[103][2]  ( .ip(n17037), .ck(clk), .q(\x[103][2] ) );
  dp_1 \x_reg[103][1]  ( .ip(n17036), .ck(clk), .q(\x[103][1] ) );
  dp_1 \x_reg[103][0]  ( .ip(n17035), .ck(clk), .q(\x[103][0] ) );
  dp_1 \x_reg[102][15]  ( .ip(n17034), .ck(clk), .q(\x[102][15] ) );
  dp_1 \x_reg[102][14]  ( .ip(n17033), .ck(clk), .q(\x[102][14] ) );
  dp_1 \x_reg[102][13]  ( .ip(n17032), .ck(clk), .q(\x[102][13] ) );
  dp_1 \x_reg[102][12]  ( .ip(n17031), .ck(clk), .q(\x[102][12] ) );
  dp_1 \x_reg[102][11]  ( .ip(n17030), .ck(clk), .q(\x[102][11] ) );
  dp_1 \x_reg[102][10]  ( .ip(n17029), .ck(clk), .q(\x[102][10] ) );
  dp_1 \x_reg[102][9]  ( .ip(n17028), .ck(clk), .q(\x[102][9] ) );
  dp_1 \x_reg[102][8]  ( .ip(n17027), .ck(clk), .q(\x[102][8] ) );
  dp_1 \x_reg[102][7]  ( .ip(n17026), .ck(clk), .q(\x[102][7] ) );
  dp_1 \x_reg[102][6]  ( .ip(n17025), .ck(clk), .q(\x[102][6] ) );
  dp_1 \x_reg[102][5]  ( .ip(n17024), .ck(clk), .q(\x[102][5] ) );
  dp_1 \x_reg[102][4]  ( .ip(n17023), .ck(clk), .q(\x[102][4] ) );
  dp_1 \x_reg[102][3]  ( .ip(n17022), .ck(clk), .q(\x[102][3] ) );
  dp_1 \x_reg[102][2]  ( .ip(n17021), .ck(clk), .q(\x[102][2] ) );
  dp_1 \x_reg[102][1]  ( .ip(n17020), .ck(clk), .q(\x[102][1] ) );
  dp_1 \x_reg[102][0]  ( .ip(n17019), .ck(clk), .q(\x[102][0] ) );
  dp_1 \x_reg[101][15]  ( .ip(n17018), .ck(clk), .q(\x[101][15] ) );
  dp_1 \x_reg[101][14]  ( .ip(n17017), .ck(clk), .q(\x[101][14] ) );
  dp_1 \x_reg[101][13]  ( .ip(n17016), .ck(clk), .q(\x[101][13] ) );
  dp_1 \x_reg[101][12]  ( .ip(n17015), .ck(clk), .q(\x[101][12] ) );
  dp_1 \x_reg[101][11]  ( .ip(n17014), .ck(clk), .q(\x[101][11] ) );
  dp_1 \x_reg[101][10]  ( .ip(n17013), .ck(clk), .q(\x[101][10] ) );
  dp_1 \x_reg[101][9]  ( .ip(n17012), .ck(clk), .q(\x[101][9] ) );
  dp_1 \x_reg[101][8]  ( .ip(n17011), .ck(clk), .q(\x[101][8] ) );
  dp_1 \x_reg[101][7]  ( .ip(n17010), .ck(clk), .q(\x[101][7] ) );
  dp_1 \x_reg[101][6]  ( .ip(n17009), .ck(clk), .q(\x[101][6] ) );
  dp_1 \x_reg[101][5]  ( .ip(n17008), .ck(clk), .q(\x[101][5] ) );
  dp_1 \x_reg[101][4]  ( .ip(n17007), .ck(clk), .q(\x[101][4] ) );
  dp_1 \x_reg[101][3]  ( .ip(n17006), .ck(clk), .q(\x[101][3] ) );
  dp_1 \x_reg[101][2]  ( .ip(n17005), .ck(clk), .q(\x[101][2] ) );
  dp_1 \x_reg[101][1]  ( .ip(n17004), .ck(clk), .q(\x[101][1] ) );
  dp_1 \x_reg[101][0]  ( .ip(n17003), .ck(clk), .q(\x[101][0] ) );
  dp_1 \x_reg[100][15]  ( .ip(n17002), .ck(clk), .q(\x[100][15] ) );
  dp_1 \x_reg[100][14]  ( .ip(n17001), .ck(clk), .q(\x[100][14] ) );
  dp_1 \x_reg[100][13]  ( .ip(n17000), .ck(clk), .q(\x[100][13] ) );
  dp_1 \x_reg[100][12]  ( .ip(n16999), .ck(clk), .q(\x[100][12] ) );
  dp_1 \x_reg[100][11]  ( .ip(n16998), .ck(clk), .q(\x[100][11] ) );
  dp_1 \x_reg[100][10]  ( .ip(n16997), .ck(clk), .q(\x[100][10] ) );
  dp_1 \x_reg[100][9]  ( .ip(n16996), .ck(clk), .q(\x[100][9] ) );
  dp_1 \x_reg[100][8]  ( .ip(n16995), .ck(clk), .q(\x[100][8] ) );
  dp_1 \x_reg[100][7]  ( .ip(n16994), .ck(clk), .q(\x[100][7] ) );
  dp_1 \x_reg[100][6]  ( .ip(n16993), .ck(clk), .q(\x[100][6] ) );
  dp_1 \x_reg[100][5]  ( .ip(n16992), .ck(clk), .q(\x[100][5] ) );
  dp_1 \x_reg[100][4]  ( .ip(n16991), .ck(clk), .q(\x[100][4] ) );
  dp_1 \x_reg[100][3]  ( .ip(n16990), .ck(clk), .q(\x[100][3] ) );
  dp_1 \x_reg[100][2]  ( .ip(n16989), .ck(clk), .q(\x[100][2] ) );
  dp_1 \x_reg[100][1]  ( .ip(n16988), .ck(clk), .q(\x[100][1] ) );
  dp_1 \x_reg[100][0]  ( .ip(n16987), .ck(clk), .q(\x[100][0] ) );
  dp_1 \x_reg[99][15]  ( .ip(n16986), .ck(clk), .q(\x[99][15] ) );
  dp_1 \x_reg[99][14]  ( .ip(n16985), .ck(clk), .q(\x[99][14] ) );
  dp_1 \x_reg[99][13]  ( .ip(n16984), .ck(clk), .q(\x[99][13] ) );
  dp_1 \x_reg[99][12]  ( .ip(n16983), .ck(clk), .q(\x[99][12] ) );
  dp_1 \x_reg[99][11]  ( .ip(n16982), .ck(clk), .q(\x[99][11] ) );
  dp_1 \x_reg[99][10]  ( .ip(n16981), .ck(clk), .q(\x[99][10] ) );
  dp_1 \x_reg[99][9]  ( .ip(n16980), .ck(clk), .q(\x[99][9] ) );
  dp_1 \x_reg[99][8]  ( .ip(n16979), .ck(clk), .q(\x[99][8] ) );
  dp_1 \x_reg[99][7]  ( .ip(n16978), .ck(clk), .q(\x[99][7] ) );
  dp_1 \x_reg[99][6]  ( .ip(n16977), .ck(clk), .q(\x[99][6] ) );
  dp_1 \x_reg[99][5]  ( .ip(n16976), .ck(clk), .q(\x[99][5] ) );
  dp_1 \x_reg[99][4]  ( .ip(n16975), .ck(clk), .q(\x[99][4] ) );
  dp_1 \x_reg[99][3]  ( .ip(n16974), .ck(clk), .q(\x[99][3] ) );
  dp_1 \x_reg[99][2]  ( .ip(n16973), .ck(clk), .q(\x[99][2] ) );
  dp_1 \x_reg[99][1]  ( .ip(n16972), .ck(clk), .q(\x[99][1] ) );
  dp_1 \x_reg[99][0]  ( .ip(n16971), .ck(clk), .q(\x[99][0] ) );
  dp_1 \x_reg[98][15]  ( .ip(n16970), .ck(clk), .q(\x[98][15] ) );
  dp_1 \x_reg[98][14]  ( .ip(n16969), .ck(clk), .q(\x[98][14] ) );
  dp_1 \x_reg[98][13]  ( .ip(n16968), .ck(clk), .q(\x[98][13] ) );
  dp_1 \x_reg[98][12]  ( .ip(n16967), .ck(clk), .q(\x[98][12] ) );
  dp_1 \x_reg[98][11]  ( .ip(n16966), .ck(clk), .q(\x[98][11] ) );
  dp_1 \x_reg[98][10]  ( .ip(n16965), .ck(clk), .q(\x[98][10] ) );
  dp_1 \x_reg[98][9]  ( .ip(n16964), .ck(clk), .q(\x[98][9] ) );
  dp_1 \x_reg[98][8]  ( .ip(n16963), .ck(clk), .q(\x[98][8] ) );
  dp_1 \x_reg[98][7]  ( .ip(n16962), .ck(clk), .q(\x[98][7] ) );
  dp_1 \x_reg[98][6]  ( .ip(n16961), .ck(clk), .q(\x[98][6] ) );
  dp_1 \x_reg[98][5]  ( .ip(n16960), .ck(clk), .q(\x[98][5] ) );
  dp_1 \x_reg[98][4]  ( .ip(n16959), .ck(clk), .q(\x[98][4] ) );
  dp_1 \x_reg[98][3]  ( .ip(n16958), .ck(clk), .q(\x[98][3] ) );
  dp_1 \x_reg[98][2]  ( .ip(n16957), .ck(clk), .q(\x[98][2] ) );
  dp_1 \x_reg[98][1]  ( .ip(n16956), .ck(clk), .q(\x[98][1] ) );
  dp_1 \x_reg[98][0]  ( .ip(n16955), .ck(clk), .q(\x[98][0] ) );
  dp_1 \x_reg[97][15]  ( .ip(n16954), .ck(clk), .q(\x[97][15] ) );
  dp_1 \x_reg[97][14]  ( .ip(n16953), .ck(clk), .q(\x[97][14] ) );
  dp_1 \x_reg[97][13]  ( .ip(n16952), .ck(clk), .q(\x[97][13] ) );
  dp_1 \x_reg[97][12]  ( .ip(n16951), .ck(clk), .q(\x[97][12] ) );
  dp_1 \x_reg[97][11]  ( .ip(n16950), .ck(clk), .q(\x[97][11] ) );
  dp_1 \x_reg[97][10]  ( .ip(n16949), .ck(clk), .q(\x[97][10] ) );
  dp_1 \x_reg[97][9]  ( .ip(n16948), .ck(clk), .q(\x[97][9] ) );
  dp_1 \x_reg[97][8]  ( .ip(n16947), .ck(clk), .q(\x[97][8] ) );
  dp_1 \x_reg[97][7]  ( .ip(n16946), .ck(clk), .q(\x[97][7] ) );
  dp_1 \x_reg[97][6]  ( .ip(n16945), .ck(clk), .q(\x[97][6] ) );
  dp_1 \x_reg[97][5]  ( .ip(n16944), .ck(clk), .q(\x[97][5] ) );
  dp_1 \x_reg[97][4]  ( .ip(n16943), .ck(clk), .q(\x[97][4] ) );
  dp_1 \x_reg[97][3]  ( .ip(n16942), .ck(clk), .q(\x[97][3] ) );
  dp_1 \x_reg[97][2]  ( .ip(n16941), .ck(clk), .q(\x[97][2] ) );
  dp_1 \x_reg[97][1]  ( .ip(n16940), .ck(clk), .q(\x[97][1] ) );
  dp_1 \x_reg[97][0]  ( .ip(n16939), .ck(clk), .q(\x[97][0] ) );
  dp_1 \x_reg[96][15]  ( .ip(n16938), .ck(clk), .q(\x[96][15] ) );
  dp_1 \x_reg[96][14]  ( .ip(n16937), .ck(clk), .q(\x[96][14] ) );
  dp_1 \x_reg[96][13]  ( .ip(n16936), .ck(clk), .q(\x[96][13] ) );
  dp_1 \x_reg[96][12]  ( .ip(n16935), .ck(clk), .q(\x[96][12] ) );
  dp_1 \x_reg[96][11]  ( .ip(n16934), .ck(clk), .q(\x[96][11] ) );
  dp_1 \x_reg[96][10]  ( .ip(n16933), .ck(clk), .q(\x[96][10] ) );
  dp_1 \x_reg[96][9]  ( .ip(n16932), .ck(clk), .q(\x[96][9] ) );
  dp_1 \x_reg[96][8]  ( .ip(n16931), .ck(clk), .q(\x[96][8] ) );
  dp_1 \x_reg[96][7]  ( .ip(n16930), .ck(clk), .q(\x[96][7] ) );
  dp_1 \x_reg[96][6]  ( .ip(n16929), .ck(clk), .q(\x[96][6] ) );
  dp_1 \x_reg[96][5]  ( .ip(n16928), .ck(clk), .q(\x[96][5] ) );
  dp_1 \x_reg[96][4]  ( .ip(n16927), .ck(clk), .q(\x[96][4] ) );
  dp_1 \x_reg[96][3]  ( .ip(n16926), .ck(clk), .q(\x[96][3] ) );
  dp_1 \x_reg[96][2]  ( .ip(n16925), .ck(clk), .q(\x[96][2] ) );
  dp_1 \x_reg[96][1]  ( .ip(n16924), .ck(clk), .q(\x[96][1] ) );
  dp_1 \x_reg[96][0]  ( .ip(n16923), .ck(clk), .q(\x[96][0] ) );
  dp_1 \x_reg[95][15]  ( .ip(n16922), .ck(clk), .q(\x[95][15] ) );
  dp_1 \x_reg[95][14]  ( .ip(n16921), .ck(clk), .q(\x[95][14] ) );
  dp_1 \x_reg[95][13]  ( .ip(n16920), .ck(clk), .q(\x[95][13] ) );
  dp_1 \x_reg[95][12]  ( .ip(n16919), .ck(clk), .q(\x[95][12] ) );
  dp_1 \x_reg[95][11]  ( .ip(n16918), .ck(clk), .q(\x[95][11] ) );
  dp_1 \x_reg[95][10]  ( .ip(n16917), .ck(clk), .q(\x[95][10] ) );
  dp_1 \x_reg[95][9]  ( .ip(n16916), .ck(clk), .q(\x[95][9] ) );
  dp_1 \x_reg[95][8]  ( .ip(n16915), .ck(clk), .q(\x[95][8] ) );
  dp_1 \x_reg[95][7]  ( .ip(n16914), .ck(clk), .q(\x[95][7] ) );
  dp_1 \x_reg[95][6]  ( .ip(n16913), .ck(clk), .q(\x[95][6] ) );
  dp_1 \x_reg[95][5]  ( .ip(n16912), .ck(clk), .q(\x[95][5] ) );
  dp_1 \x_reg[95][4]  ( .ip(n16911), .ck(clk), .q(\x[95][4] ) );
  dp_1 \x_reg[95][3]  ( .ip(n16910), .ck(clk), .q(\x[95][3] ) );
  dp_1 \x_reg[95][2]  ( .ip(n16909), .ck(clk), .q(\x[95][2] ) );
  dp_1 \x_reg[95][1]  ( .ip(n16908), .ck(clk), .q(\x[95][1] ) );
  dp_1 \x_reg[95][0]  ( .ip(n16907), .ck(clk), .q(\x[95][0] ) );
  dp_1 \x_reg[94][15]  ( .ip(n16906), .ck(clk), .q(\x[94][15] ) );
  dp_1 \x_reg[94][14]  ( .ip(n16905), .ck(clk), .q(\x[94][14] ) );
  dp_1 \x_reg[94][13]  ( .ip(n16904), .ck(clk), .q(\x[94][13] ) );
  dp_1 \x_reg[94][12]  ( .ip(n16903), .ck(clk), .q(\x[94][12] ) );
  dp_1 \x_reg[94][11]  ( .ip(n16902), .ck(clk), .q(\x[94][11] ) );
  dp_1 \x_reg[94][10]  ( .ip(n16901), .ck(clk), .q(\x[94][10] ) );
  dp_1 \x_reg[94][9]  ( .ip(n16900), .ck(clk), .q(\x[94][9] ) );
  dp_1 \x_reg[94][8]  ( .ip(n16899), .ck(clk), .q(\x[94][8] ) );
  dp_1 \x_reg[94][7]  ( .ip(n16898), .ck(clk), .q(\x[94][7] ) );
  dp_1 \x_reg[94][6]  ( .ip(n16897), .ck(clk), .q(\x[94][6] ) );
  dp_1 \x_reg[94][5]  ( .ip(n16896), .ck(clk), .q(\x[94][5] ) );
  dp_1 \x_reg[94][4]  ( .ip(n16895), .ck(clk), .q(\x[94][4] ) );
  dp_1 \x_reg[94][3]  ( .ip(n16894), .ck(clk), .q(\x[94][3] ) );
  dp_1 \x_reg[94][2]  ( .ip(n16893), .ck(clk), .q(\x[94][2] ) );
  dp_1 \x_reg[94][1]  ( .ip(n16892), .ck(clk), .q(\x[94][1] ) );
  dp_1 \x_reg[94][0]  ( .ip(n16891), .ck(clk), .q(\x[94][0] ) );
  dp_1 \x_reg[93][15]  ( .ip(n16890), .ck(clk), .q(\x[93][15] ) );
  dp_1 \x_reg[93][14]  ( .ip(n16889), .ck(clk), .q(\x[93][14] ) );
  dp_1 \x_reg[93][13]  ( .ip(n16888), .ck(clk), .q(\x[93][13] ) );
  dp_1 \x_reg[93][12]  ( .ip(n16887), .ck(clk), .q(\x[93][12] ) );
  dp_1 \x_reg[93][11]  ( .ip(n16886), .ck(clk), .q(\x[93][11] ) );
  dp_1 \x_reg[93][10]  ( .ip(n16885), .ck(clk), .q(\x[93][10] ) );
  dp_1 \x_reg[93][9]  ( .ip(n16884), .ck(clk), .q(\x[93][9] ) );
  dp_1 \x_reg[93][8]  ( .ip(n16883), .ck(clk), .q(\x[93][8] ) );
  dp_1 \x_reg[93][7]  ( .ip(n16882), .ck(clk), .q(\x[93][7] ) );
  dp_1 \x_reg[93][6]  ( .ip(n16881), .ck(clk), .q(\x[93][6] ) );
  dp_1 \x_reg[93][5]  ( .ip(n16880), .ck(clk), .q(\x[93][5] ) );
  dp_1 \x_reg[93][4]  ( .ip(n16879), .ck(clk), .q(\x[93][4] ) );
  dp_1 \x_reg[93][3]  ( .ip(n16878), .ck(clk), .q(\x[93][3] ) );
  dp_1 \x_reg[93][2]  ( .ip(n16877), .ck(clk), .q(\x[93][2] ) );
  dp_1 \x_reg[93][1]  ( .ip(n16876), .ck(clk), .q(\x[93][1] ) );
  dp_1 \x_reg[93][0]  ( .ip(n16875), .ck(clk), .q(\x[93][0] ) );
  dp_1 \x_reg[92][15]  ( .ip(n16874), .ck(clk), .q(\x[92][15] ) );
  dp_1 \x_reg[92][14]  ( .ip(n16873), .ck(clk), .q(\x[92][14] ) );
  dp_1 \x_reg[92][13]  ( .ip(n16872), .ck(clk), .q(\x[92][13] ) );
  dp_1 \x_reg[92][12]  ( .ip(n16871), .ck(clk), .q(\x[92][12] ) );
  dp_1 \x_reg[92][11]  ( .ip(n16870), .ck(clk), .q(\x[92][11] ) );
  dp_1 \x_reg[92][10]  ( .ip(n16869), .ck(clk), .q(\x[92][10] ) );
  dp_1 \x_reg[92][9]  ( .ip(n16868), .ck(clk), .q(\x[92][9] ) );
  dp_1 \x_reg[92][8]  ( .ip(n16867), .ck(clk), .q(\x[92][8] ) );
  dp_1 \x_reg[92][7]  ( .ip(n16866), .ck(clk), .q(\x[92][7] ) );
  dp_1 \x_reg[92][6]  ( .ip(n16865), .ck(clk), .q(\x[92][6] ) );
  dp_1 \x_reg[92][5]  ( .ip(n16864), .ck(clk), .q(\x[92][5] ) );
  dp_1 \x_reg[92][4]  ( .ip(n16863), .ck(clk), .q(\x[92][4] ) );
  dp_1 \x_reg[92][3]  ( .ip(n16862), .ck(clk), .q(\x[92][3] ) );
  dp_1 \x_reg[92][2]  ( .ip(n16861), .ck(clk), .q(\x[92][2] ) );
  dp_1 \x_reg[92][1]  ( .ip(n16860), .ck(clk), .q(\x[92][1] ) );
  dp_1 \x_reg[92][0]  ( .ip(n16859), .ck(clk), .q(\x[92][0] ) );
  dp_1 \x_reg[91][15]  ( .ip(n16858), .ck(clk), .q(\x[91][15] ) );
  dp_1 \x_reg[91][14]  ( .ip(n16857), .ck(clk), .q(\x[91][14] ) );
  dp_1 \x_reg[91][13]  ( .ip(n16856), .ck(clk), .q(\x[91][13] ) );
  dp_1 \x_reg[91][12]  ( .ip(n16855), .ck(clk), .q(\x[91][12] ) );
  dp_1 \x_reg[91][11]  ( .ip(n16854), .ck(clk), .q(\x[91][11] ) );
  dp_1 \x_reg[91][10]  ( .ip(n16853), .ck(clk), .q(\x[91][10] ) );
  dp_1 \x_reg[91][9]  ( .ip(n16852), .ck(clk), .q(\x[91][9] ) );
  dp_1 \x_reg[91][8]  ( .ip(n16851), .ck(clk), .q(\x[91][8] ) );
  dp_1 \x_reg[91][7]  ( .ip(n16850), .ck(clk), .q(\x[91][7] ) );
  dp_1 \x_reg[91][6]  ( .ip(n16849), .ck(clk), .q(\x[91][6] ) );
  dp_1 \x_reg[91][5]  ( .ip(n16848), .ck(clk), .q(\x[91][5] ) );
  dp_1 \x_reg[91][4]  ( .ip(n16847), .ck(clk), .q(\x[91][4] ) );
  dp_1 \x_reg[91][3]  ( .ip(n16846), .ck(clk), .q(\x[91][3] ) );
  dp_1 \x_reg[91][2]  ( .ip(n16845), .ck(clk), .q(\x[91][2] ) );
  dp_1 \x_reg[91][1]  ( .ip(n16844), .ck(clk), .q(\x[91][1] ) );
  dp_1 \x_reg[91][0]  ( .ip(n16843), .ck(clk), .q(\x[91][0] ) );
  dp_1 \x_reg[90][15]  ( .ip(n16842), .ck(clk), .q(\x[90][15] ) );
  dp_1 \x_reg[90][14]  ( .ip(n16841), .ck(clk), .q(\x[90][14] ) );
  dp_1 \x_reg[90][13]  ( .ip(n16840), .ck(clk), .q(\x[90][13] ) );
  dp_1 \x_reg[90][12]  ( .ip(n16839), .ck(clk), .q(\x[90][12] ) );
  dp_1 \x_reg[90][11]  ( .ip(n16838), .ck(clk), .q(\x[90][11] ) );
  dp_1 \x_reg[90][10]  ( .ip(n16837), .ck(clk), .q(\x[90][10] ) );
  dp_1 \x_reg[90][9]  ( .ip(n16836), .ck(clk), .q(\x[90][9] ) );
  dp_1 \x_reg[90][8]  ( .ip(n16835), .ck(clk), .q(\x[90][8] ) );
  dp_1 \x_reg[90][7]  ( .ip(n16834), .ck(clk), .q(\x[90][7] ) );
  dp_1 \x_reg[90][6]  ( .ip(n16833), .ck(clk), .q(\x[90][6] ) );
  dp_1 \x_reg[90][5]  ( .ip(n16832), .ck(clk), .q(\x[90][5] ) );
  dp_1 \x_reg[90][4]  ( .ip(n16831), .ck(clk), .q(\x[90][4] ) );
  dp_1 \x_reg[90][3]  ( .ip(n16830), .ck(clk), .q(\x[90][3] ) );
  dp_1 \x_reg[90][2]  ( .ip(n16829), .ck(clk), .q(\x[90][2] ) );
  dp_1 \x_reg[90][1]  ( .ip(n16828), .ck(clk), .q(\x[90][1] ) );
  dp_1 \x_reg[90][0]  ( .ip(n16827), .ck(clk), .q(\x[90][0] ) );
  dp_1 \x_reg[89][15]  ( .ip(n16826), .ck(clk), .q(\x[89][15] ) );
  dp_1 \x_reg[89][14]  ( .ip(n16825), .ck(clk), .q(\x[89][14] ) );
  dp_1 \x_reg[89][13]  ( .ip(n16824), .ck(clk), .q(\x[89][13] ) );
  dp_1 \x_reg[89][12]  ( .ip(n16823), .ck(clk), .q(\x[89][12] ) );
  dp_1 \x_reg[89][11]  ( .ip(n16822), .ck(clk), .q(\x[89][11] ) );
  dp_1 \x_reg[89][10]  ( .ip(n16821), .ck(clk), .q(\x[89][10] ) );
  dp_1 \x_reg[89][9]  ( .ip(n16820), .ck(clk), .q(\x[89][9] ) );
  dp_1 \x_reg[89][8]  ( .ip(n16819), .ck(clk), .q(\x[89][8] ) );
  dp_1 \x_reg[89][7]  ( .ip(n16818), .ck(clk), .q(\x[89][7] ) );
  dp_1 \x_reg[89][6]  ( .ip(n16817), .ck(clk), .q(\x[89][6] ) );
  dp_1 \x_reg[89][5]  ( .ip(n16816), .ck(clk), .q(\x[89][5] ) );
  dp_1 \x_reg[89][4]  ( .ip(n16815), .ck(clk), .q(\x[89][4] ) );
  dp_1 \x_reg[89][3]  ( .ip(n16814), .ck(clk), .q(\x[89][3] ) );
  dp_1 \x_reg[89][2]  ( .ip(n16813), .ck(clk), .q(\x[89][2] ) );
  dp_1 \x_reg[89][1]  ( .ip(n16812), .ck(clk), .q(\x[89][1] ) );
  dp_1 \x_reg[89][0]  ( .ip(n16811), .ck(clk), .q(\x[89][0] ) );
  dp_1 \x_reg[88][15]  ( .ip(n16810), .ck(clk), .q(\x[88][15] ) );
  dp_1 \x_reg[88][14]  ( .ip(n16809), .ck(clk), .q(\x[88][14] ) );
  dp_1 \x_reg[88][13]  ( .ip(n16808), .ck(clk), .q(\x[88][13] ) );
  dp_1 \x_reg[88][12]  ( .ip(n16807), .ck(clk), .q(\x[88][12] ) );
  dp_1 \x_reg[88][11]  ( .ip(n16806), .ck(clk), .q(\x[88][11] ) );
  dp_1 \x_reg[88][10]  ( .ip(n16805), .ck(clk), .q(\x[88][10] ) );
  dp_1 \x_reg[88][9]  ( .ip(n16804), .ck(clk), .q(\x[88][9] ) );
  dp_1 \x_reg[88][8]  ( .ip(n16803), .ck(clk), .q(\x[88][8] ) );
  dp_1 \x_reg[88][7]  ( .ip(n16802), .ck(clk), .q(\x[88][7] ) );
  dp_1 \x_reg[88][6]  ( .ip(n16801), .ck(clk), .q(\x[88][6] ) );
  dp_1 \x_reg[88][5]  ( .ip(n16800), .ck(clk), .q(\x[88][5] ) );
  dp_1 \x_reg[88][4]  ( .ip(n16799), .ck(clk), .q(\x[88][4] ) );
  dp_1 \x_reg[88][3]  ( .ip(n16798), .ck(clk), .q(\x[88][3] ) );
  dp_1 \x_reg[88][2]  ( .ip(n16797), .ck(clk), .q(\x[88][2] ) );
  dp_1 \x_reg[88][1]  ( .ip(n16796), .ck(clk), .q(\x[88][1] ) );
  dp_1 \x_reg[88][0]  ( .ip(n16795), .ck(clk), .q(\x[88][0] ) );
  dp_1 \x_reg[87][15]  ( .ip(n16794), .ck(clk), .q(\x[87][15] ) );
  dp_1 \x_reg[87][14]  ( .ip(n16793), .ck(clk), .q(\x[87][14] ) );
  dp_1 \x_reg[87][13]  ( .ip(n16792), .ck(clk), .q(\x[87][13] ) );
  dp_1 \x_reg[87][12]  ( .ip(n16791), .ck(clk), .q(\x[87][12] ) );
  dp_1 \x_reg[87][11]  ( .ip(n16790), .ck(clk), .q(\x[87][11] ) );
  dp_1 \x_reg[87][10]  ( .ip(n16789), .ck(clk), .q(\x[87][10] ) );
  dp_1 \x_reg[87][9]  ( .ip(n16788), .ck(clk), .q(\x[87][9] ) );
  dp_1 \x_reg[87][8]  ( .ip(n16787), .ck(clk), .q(\x[87][8] ) );
  dp_1 \x_reg[87][7]  ( .ip(n16786), .ck(clk), .q(\x[87][7] ) );
  dp_1 \x_reg[87][6]  ( .ip(n16785), .ck(clk), .q(\x[87][6] ) );
  dp_1 \x_reg[87][5]  ( .ip(n16784), .ck(clk), .q(\x[87][5] ) );
  dp_1 \x_reg[87][4]  ( .ip(n16783), .ck(clk), .q(\x[87][4] ) );
  dp_1 \x_reg[87][3]  ( .ip(n16782), .ck(clk), .q(\x[87][3] ) );
  dp_1 \x_reg[87][2]  ( .ip(n16781), .ck(clk), .q(\x[87][2] ) );
  dp_1 \x_reg[87][1]  ( .ip(n16780), .ck(clk), .q(\x[87][1] ) );
  dp_1 \x_reg[87][0]  ( .ip(n16779), .ck(clk), .q(\x[87][0] ) );
  dp_1 \x_reg[86][15]  ( .ip(n16778), .ck(clk), .q(\x[86][15] ) );
  dp_1 \x_reg[86][14]  ( .ip(n16777), .ck(clk), .q(\x[86][14] ) );
  dp_1 \x_reg[86][13]  ( .ip(n16776), .ck(clk), .q(\x[86][13] ) );
  dp_1 \x_reg[86][12]  ( .ip(n16775), .ck(clk), .q(\x[86][12] ) );
  dp_1 \x_reg[86][11]  ( .ip(n16774), .ck(clk), .q(\x[86][11] ) );
  dp_1 \x_reg[86][10]  ( .ip(n16773), .ck(clk), .q(\x[86][10] ) );
  dp_1 \x_reg[86][9]  ( .ip(n16772), .ck(clk), .q(\x[86][9] ) );
  dp_1 \x_reg[86][8]  ( .ip(n16771), .ck(clk), .q(\x[86][8] ) );
  dp_1 \x_reg[86][7]  ( .ip(n16770), .ck(clk), .q(\x[86][7] ) );
  dp_1 \x_reg[86][6]  ( .ip(n16769), .ck(clk), .q(\x[86][6] ) );
  dp_1 \x_reg[86][5]  ( .ip(n16768), .ck(clk), .q(\x[86][5] ) );
  dp_1 \x_reg[86][4]  ( .ip(n16767), .ck(clk), .q(\x[86][4] ) );
  dp_1 \x_reg[86][3]  ( .ip(n16766), .ck(clk), .q(\x[86][3] ) );
  dp_1 \x_reg[86][2]  ( .ip(n16765), .ck(clk), .q(\x[86][2] ) );
  dp_1 \x_reg[86][1]  ( .ip(n16764), .ck(clk), .q(\x[86][1] ) );
  dp_1 \x_reg[86][0]  ( .ip(n16763), .ck(clk), .q(\x[86][0] ) );
  dp_1 \x_reg[85][15]  ( .ip(n16762), .ck(clk), .q(\x[85][15] ) );
  dp_1 \x_reg[85][14]  ( .ip(n16761), .ck(clk), .q(\x[85][14] ) );
  dp_1 \x_reg[85][13]  ( .ip(n16760), .ck(clk), .q(\x[85][13] ) );
  dp_1 \x_reg[85][12]  ( .ip(n16759), .ck(clk), .q(\x[85][12] ) );
  dp_1 \x_reg[85][11]  ( .ip(n16758), .ck(clk), .q(\x[85][11] ) );
  dp_1 \x_reg[85][10]  ( .ip(n16757), .ck(clk), .q(\x[85][10] ) );
  dp_1 \x_reg[85][9]  ( .ip(n16756), .ck(clk), .q(\x[85][9] ) );
  dp_1 \x_reg[85][8]  ( .ip(n16755), .ck(clk), .q(\x[85][8] ) );
  dp_1 \x_reg[85][7]  ( .ip(n16754), .ck(clk), .q(\x[85][7] ) );
  dp_1 \x_reg[85][6]  ( .ip(n16753), .ck(clk), .q(\x[85][6] ) );
  dp_1 \x_reg[85][5]  ( .ip(n16752), .ck(clk), .q(\x[85][5] ) );
  dp_1 \x_reg[85][4]  ( .ip(n16751), .ck(clk), .q(\x[85][4] ) );
  dp_1 \x_reg[85][3]  ( .ip(n16750), .ck(clk), .q(\x[85][3] ) );
  dp_1 \x_reg[85][2]  ( .ip(n16749), .ck(clk), .q(\x[85][2] ) );
  dp_1 \x_reg[85][1]  ( .ip(n16748), .ck(clk), .q(\x[85][1] ) );
  dp_1 \x_reg[85][0]  ( .ip(n16747), .ck(clk), .q(\x[85][0] ) );
  dp_1 \x_reg[84][15]  ( .ip(n16746), .ck(clk), .q(\x[84][15] ) );
  dp_1 \x_reg[84][14]  ( .ip(n16745), .ck(clk), .q(\x[84][14] ) );
  dp_1 \x_reg[84][13]  ( .ip(n16744), .ck(clk), .q(\x[84][13] ) );
  dp_1 \x_reg[84][12]  ( .ip(n16743), .ck(clk), .q(\x[84][12] ) );
  dp_1 \x_reg[84][11]  ( .ip(n16742), .ck(clk), .q(\x[84][11] ) );
  dp_1 \x_reg[84][10]  ( .ip(n16741), .ck(clk), .q(\x[84][10] ) );
  dp_1 \x_reg[84][9]  ( .ip(n16740), .ck(clk), .q(\x[84][9] ) );
  dp_1 \x_reg[84][8]  ( .ip(n16739), .ck(clk), .q(\x[84][8] ) );
  dp_1 \x_reg[84][7]  ( .ip(n16738), .ck(clk), .q(\x[84][7] ) );
  dp_1 \x_reg[84][6]  ( .ip(n16737), .ck(clk), .q(\x[84][6] ) );
  dp_1 \x_reg[84][5]  ( .ip(n16736), .ck(clk), .q(\x[84][5] ) );
  dp_1 \x_reg[84][4]  ( .ip(n16735), .ck(clk), .q(\x[84][4] ) );
  dp_1 \x_reg[84][3]  ( .ip(n16734), .ck(clk), .q(\x[84][3] ) );
  dp_1 \x_reg[84][2]  ( .ip(n16733), .ck(clk), .q(\x[84][2] ) );
  dp_1 \x_reg[84][1]  ( .ip(n16732), .ck(clk), .q(\x[84][1] ) );
  dp_1 \x_reg[84][0]  ( .ip(n16731), .ck(clk), .q(\x[84][0] ) );
  dp_1 \x_reg[83][15]  ( .ip(n16730), .ck(clk), .q(\x[83][15] ) );
  dp_1 \x_reg[83][14]  ( .ip(n16729), .ck(clk), .q(\x[83][14] ) );
  dp_1 \x_reg[83][13]  ( .ip(n16728), .ck(clk), .q(\x[83][13] ) );
  dp_1 \x_reg[83][12]  ( .ip(n16727), .ck(clk), .q(\x[83][12] ) );
  dp_1 \x_reg[83][11]  ( .ip(n16726), .ck(clk), .q(\x[83][11] ) );
  dp_1 \x_reg[83][10]  ( .ip(n16725), .ck(clk), .q(\x[83][10] ) );
  dp_1 \x_reg[83][9]  ( .ip(n16724), .ck(clk), .q(\x[83][9] ) );
  dp_1 \x_reg[83][8]  ( .ip(n16723), .ck(clk), .q(\x[83][8] ) );
  dp_1 \x_reg[83][7]  ( .ip(n16722), .ck(clk), .q(\x[83][7] ) );
  dp_1 \x_reg[83][6]  ( .ip(n16721), .ck(clk), .q(\x[83][6] ) );
  dp_1 \x_reg[83][5]  ( .ip(n16720), .ck(clk), .q(\x[83][5] ) );
  dp_1 \x_reg[83][4]  ( .ip(n16719), .ck(clk), .q(\x[83][4] ) );
  dp_1 \x_reg[83][3]  ( .ip(n16718), .ck(clk), .q(\x[83][3] ) );
  dp_1 \x_reg[83][2]  ( .ip(n16717), .ck(clk), .q(\x[83][2] ) );
  dp_1 \x_reg[83][1]  ( .ip(n16716), .ck(clk), .q(\x[83][1] ) );
  dp_1 \x_reg[83][0]  ( .ip(n16715), .ck(clk), .q(\x[83][0] ) );
  dp_1 \x_reg[82][15]  ( .ip(n16714), .ck(clk), .q(\x[82][15] ) );
  dp_1 \x_reg[82][14]  ( .ip(n16713), .ck(clk), .q(\x[82][14] ) );
  dp_1 \x_reg[82][13]  ( .ip(n16712), .ck(clk), .q(\x[82][13] ) );
  dp_1 \x_reg[82][12]  ( .ip(n16711), .ck(clk), .q(\x[82][12] ) );
  dp_1 \x_reg[82][11]  ( .ip(n16710), .ck(clk), .q(\x[82][11] ) );
  dp_1 \x_reg[82][10]  ( .ip(n16709), .ck(clk), .q(\x[82][10] ) );
  dp_1 \x_reg[82][9]  ( .ip(n16708), .ck(clk), .q(\x[82][9] ) );
  dp_1 \x_reg[82][8]  ( .ip(n16707), .ck(clk), .q(\x[82][8] ) );
  dp_1 \x_reg[82][7]  ( .ip(n16706), .ck(clk), .q(\x[82][7] ) );
  dp_1 \x_reg[82][6]  ( .ip(n16705), .ck(clk), .q(\x[82][6] ) );
  dp_1 \x_reg[82][5]  ( .ip(n16704), .ck(clk), .q(\x[82][5] ) );
  dp_1 \x_reg[82][4]  ( .ip(n16703), .ck(clk), .q(\x[82][4] ) );
  dp_1 \x_reg[82][3]  ( .ip(n16702), .ck(clk), .q(\x[82][3] ) );
  dp_1 \x_reg[82][2]  ( .ip(n16701), .ck(clk), .q(\x[82][2] ) );
  dp_1 \x_reg[82][1]  ( .ip(n16700), .ck(clk), .q(\x[82][1] ) );
  dp_1 \x_reg[82][0]  ( .ip(n16699), .ck(clk), .q(\x[82][0] ) );
  dp_1 \x_reg[81][15]  ( .ip(n16698), .ck(clk), .q(\x[81][15] ) );
  dp_1 \x_reg[81][14]  ( .ip(n16697), .ck(clk), .q(\x[81][14] ) );
  dp_1 \x_reg[81][13]  ( .ip(n16696), .ck(clk), .q(\x[81][13] ) );
  dp_1 \x_reg[81][12]  ( .ip(n16695), .ck(clk), .q(\x[81][12] ) );
  dp_1 \x_reg[81][11]  ( .ip(n16694), .ck(clk), .q(\x[81][11] ) );
  dp_1 \x_reg[81][10]  ( .ip(n16693), .ck(clk), .q(\x[81][10] ) );
  dp_1 \x_reg[81][9]  ( .ip(n16692), .ck(clk), .q(\x[81][9] ) );
  dp_1 \x_reg[81][8]  ( .ip(n16691), .ck(clk), .q(\x[81][8] ) );
  dp_1 \x_reg[81][7]  ( .ip(n16690), .ck(clk), .q(\x[81][7] ) );
  dp_1 \x_reg[81][6]  ( .ip(n16689), .ck(clk), .q(\x[81][6] ) );
  dp_1 \x_reg[81][5]  ( .ip(n16688), .ck(clk), .q(\x[81][5] ) );
  dp_1 \x_reg[81][4]  ( .ip(n16687), .ck(clk), .q(\x[81][4] ) );
  dp_1 \x_reg[81][3]  ( .ip(n16686), .ck(clk), .q(\x[81][3] ) );
  dp_1 \x_reg[81][2]  ( .ip(n16685), .ck(clk), .q(\x[81][2] ) );
  dp_1 \x_reg[81][1]  ( .ip(n16684), .ck(clk), .q(\x[81][1] ) );
  dp_1 \x_reg[81][0]  ( .ip(n16683), .ck(clk), .q(\x[81][0] ) );
  dp_1 \x_reg[80][15]  ( .ip(n16682), .ck(clk), .q(\x[80][15] ) );
  dp_1 \x_reg[80][14]  ( .ip(n16681), .ck(clk), .q(\x[80][14] ) );
  dp_1 \x_reg[80][13]  ( .ip(n16680), .ck(clk), .q(\x[80][13] ) );
  dp_1 \x_reg[80][12]  ( .ip(n16679), .ck(clk), .q(\x[80][12] ) );
  dp_1 \x_reg[80][11]  ( .ip(n16678), .ck(clk), .q(\x[80][11] ) );
  dp_1 \x_reg[80][10]  ( .ip(n16677), .ck(clk), .q(\x[80][10] ) );
  dp_1 \x_reg[80][9]  ( .ip(n16676), .ck(clk), .q(\x[80][9] ) );
  dp_1 \x_reg[80][8]  ( .ip(n16675), .ck(clk), .q(\x[80][8] ) );
  dp_1 \x_reg[80][7]  ( .ip(n16674), .ck(clk), .q(\x[80][7] ) );
  dp_1 \x_reg[80][6]  ( .ip(n16673), .ck(clk), .q(\x[80][6] ) );
  dp_1 \x_reg[80][5]  ( .ip(n16672), .ck(clk), .q(\x[80][5] ) );
  dp_1 \x_reg[80][4]  ( .ip(n16671), .ck(clk), .q(\x[80][4] ) );
  dp_1 \x_reg[80][3]  ( .ip(n16670), .ck(clk), .q(\x[80][3] ) );
  dp_1 \x_reg[80][2]  ( .ip(n16669), .ck(clk), .q(\x[80][2] ) );
  dp_1 \x_reg[80][1]  ( .ip(n16668), .ck(clk), .q(\x[80][1] ) );
  dp_1 \x_reg[80][0]  ( .ip(n16667), .ck(clk), .q(\x[80][0] ) );
  dp_1 \x_reg[79][15]  ( .ip(n16666), .ck(clk), .q(\x[79][15] ) );
  dp_1 \x_reg[79][14]  ( .ip(n16665), .ck(clk), .q(\x[79][14] ) );
  dp_1 \x_reg[79][13]  ( .ip(n16664), .ck(clk), .q(\x[79][13] ) );
  dp_1 \x_reg[79][12]  ( .ip(n16663), .ck(clk), .q(\x[79][12] ) );
  dp_1 \x_reg[79][11]  ( .ip(n16662), .ck(clk), .q(\x[79][11] ) );
  dp_1 \x_reg[79][10]  ( .ip(n16661), .ck(clk), .q(\x[79][10] ) );
  dp_1 \x_reg[79][9]  ( .ip(n16660), .ck(clk), .q(\x[79][9] ) );
  dp_1 \x_reg[79][8]  ( .ip(n16659), .ck(clk), .q(\x[79][8] ) );
  dp_1 \x_reg[79][7]  ( .ip(n16658), .ck(clk), .q(\x[79][7] ) );
  dp_1 \x_reg[79][6]  ( .ip(n16657), .ck(clk), .q(\x[79][6] ) );
  dp_1 \x_reg[79][5]  ( .ip(n16656), .ck(clk), .q(\x[79][5] ) );
  dp_1 \x_reg[79][4]  ( .ip(n16655), .ck(clk), .q(\x[79][4] ) );
  dp_1 \x_reg[79][3]  ( .ip(n16654), .ck(clk), .q(\x[79][3] ) );
  dp_1 \x_reg[79][2]  ( .ip(n16653), .ck(clk), .q(\x[79][2] ) );
  dp_1 \x_reg[79][1]  ( .ip(n16652), .ck(clk), .q(\x[79][1] ) );
  dp_1 \x_reg[79][0]  ( .ip(n16651), .ck(clk), .q(\x[79][0] ) );
  dp_1 \x_reg[78][15]  ( .ip(n16650), .ck(clk), .q(\x[78][15] ) );
  dp_1 \x_reg[78][14]  ( .ip(n16649), .ck(clk), .q(\x[78][14] ) );
  dp_1 \x_reg[78][13]  ( .ip(n16648), .ck(clk), .q(\x[78][13] ) );
  dp_1 \x_reg[78][12]  ( .ip(n16647), .ck(clk), .q(\x[78][12] ) );
  dp_1 \x_reg[78][11]  ( .ip(n16646), .ck(clk), .q(\x[78][11] ) );
  dp_1 \x_reg[78][10]  ( .ip(n16645), .ck(clk), .q(\x[78][10] ) );
  dp_1 \x_reg[78][9]  ( .ip(n16644), .ck(clk), .q(\x[78][9] ) );
  dp_1 \x_reg[78][8]  ( .ip(n16643), .ck(clk), .q(\x[78][8] ) );
  dp_1 \x_reg[78][7]  ( .ip(n16642), .ck(clk), .q(\x[78][7] ) );
  dp_1 \x_reg[78][6]  ( .ip(n16641), .ck(clk), .q(\x[78][6] ) );
  dp_1 \x_reg[78][5]  ( .ip(n16640), .ck(clk), .q(\x[78][5] ) );
  dp_1 \x_reg[78][4]  ( .ip(n16639), .ck(clk), .q(\x[78][4] ) );
  dp_1 \x_reg[78][3]  ( .ip(n16638), .ck(clk), .q(\x[78][3] ) );
  dp_1 \x_reg[78][2]  ( .ip(n16637), .ck(clk), .q(\x[78][2] ) );
  dp_1 \x_reg[78][1]  ( .ip(n16636), .ck(clk), .q(\x[78][1] ) );
  dp_1 \x_reg[78][0]  ( .ip(n16635), .ck(clk), .q(\x[78][0] ) );
  dp_1 \x_reg[77][15]  ( .ip(n16634), .ck(clk), .q(\x[77][15] ) );
  dp_1 \x_reg[77][14]  ( .ip(n16633), .ck(clk), .q(\x[77][14] ) );
  dp_1 \x_reg[77][13]  ( .ip(n16632), .ck(clk), .q(\x[77][13] ) );
  dp_1 \x_reg[77][12]  ( .ip(n16631), .ck(clk), .q(\x[77][12] ) );
  dp_1 \x_reg[77][11]  ( .ip(n16630), .ck(clk), .q(\x[77][11] ) );
  dp_1 \x_reg[77][10]  ( .ip(n16629), .ck(clk), .q(\x[77][10] ) );
  dp_1 \x_reg[77][9]  ( .ip(n16628), .ck(clk), .q(\x[77][9] ) );
  dp_1 \x_reg[77][8]  ( .ip(n16627), .ck(clk), .q(\x[77][8] ) );
  dp_1 \x_reg[77][7]  ( .ip(n16626), .ck(clk), .q(\x[77][7] ) );
  dp_1 \x_reg[77][6]  ( .ip(n16625), .ck(clk), .q(\x[77][6] ) );
  dp_1 \x_reg[77][5]  ( .ip(n16624), .ck(clk), .q(\x[77][5] ) );
  dp_1 \x_reg[77][4]  ( .ip(n16623), .ck(clk), .q(\x[77][4] ) );
  dp_1 \x_reg[77][3]  ( .ip(n16622), .ck(clk), .q(\x[77][3] ) );
  dp_1 \x_reg[77][2]  ( .ip(n16621), .ck(clk), .q(\x[77][2] ) );
  dp_1 \x_reg[77][1]  ( .ip(n16620), .ck(clk), .q(\x[77][1] ) );
  dp_1 \x_reg[77][0]  ( .ip(n16619), .ck(clk), .q(\x[77][0] ) );
  dp_1 \x_reg[76][15]  ( .ip(n16618), .ck(clk), .q(\x[76][15] ) );
  dp_1 \x_reg[76][14]  ( .ip(n16617), .ck(clk), .q(\x[76][14] ) );
  dp_1 \x_reg[76][13]  ( .ip(n16616), .ck(clk), .q(\x[76][13] ) );
  dp_1 \x_reg[76][12]  ( .ip(n16615), .ck(clk), .q(\x[76][12] ) );
  dp_1 \x_reg[76][11]  ( .ip(n16614), .ck(clk), .q(\x[76][11] ) );
  dp_1 \x_reg[76][10]  ( .ip(n16613), .ck(clk), .q(\x[76][10] ) );
  dp_1 \x_reg[76][9]  ( .ip(n16612), .ck(clk), .q(\x[76][9] ) );
  dp_1 \x_reg[76][8]  ( .ip(n16611), .ck(clk), .q(\x[76][8] ) );
  dp_1 \x_reg[76][7]  ( .ip(n16610), .ck(clk), .q(\x[76][7] ) );
  dp_1 \x_reg[76][6]  ( .ip(n16609), .ck(clk), .q(\x[76][6] ) );
  dp_1 \x_reg[76][5]  ( .ip(n16608), .ck(clk), .q(\x[76][5] ) );
  dp_1 \x_reg[76][4]  ( .ip(n16607), .ck(clk), .q(\x[76][4] ) );
  dp_1 \x_reg[76][3]  ( .ip(n16606), .ck(clk), .q(\x[76][3] ) );
  dp_1 \x_reg[76][2]  ( .ip(n16605), .ck(clk), .q(\x[76][2] ) );
  dp_1 \x_reg[76][1]  ( .ip(n16604), .ck(clk), .q(\x[76][1] ) );
  dp_1 \x_reg[76][0]  ( .ip(n16603), .ck(clk), .q(\x[76][0] ) );
  dp_1 \x_reg[75][15]  ( .ip(n16602), .ck(clk), .q(\x[75][15] ) );
  dp_1 \x_reg[75][14]  ( .ip(n16601), .ck(clk), .q(\x[75][14] ) );
  dp_1 \x_reg[75][13]  ( .ip(n16600), .ck(clk), .q(\x[75][13] ) );
  dp_1 \x_reg[75][12]  ( .ip(n16599), .ck(clk), .q(\x[75][12] ) );
  dp_1 \x_reg[75][11]  ( .ip(n16598), .ck(clk), .q(\x[75][11] ) );
  dp_1 \x_reg[75][10]  ( .ip(n16597), .ck(clk), .q(\x[75][10] ) );
  dp_1 \x_reg[75][9]  ( .ip(n16596), .ck(clk), .q(\x[75][9] ) );
  dp_1 \x_reg[75][8]  ( .ip(n16595), .ck(clk), .q(\x[75][8] ) );
  dp_1 \x_reg[75][7]  ( .ip(n16594), .ck(clk), .q(\x[75][7] ) );
  dp_1 \x_reg[75][6]  ( .ip(n16593), .ck(clk), .q(\x[75][6] ) );
  dp_1 \x_reg[75][5]  ( .ip(n16592), .ck(clk), .q(\x[75][5] ) );
  dp_1 \x_reg[75][4]  ( .ip(n16591), .ck(clk), .q(\x[75][4] ) );
  dp_1 \x_reg[75][3]  ( .ip(n16590), .ck(clk), .q(\x[75][3] ) );
  dp_1 \x_reg[75][2]  ( .ip(n16589), .ck(clk), .q(\x[75][2] ) );
  dp_1 \x_reg[75][1]  ( .ip(n16588), .ck(clk), .q(\x[75][1] ) );
  dp_1 \x_reg[75][0]  ( .ip(n16587), .ck(clk), .q(\x[75][0] ) );
  dp_1 \x_reg[74][15]  ( .ip(n16586), .ck(clk), .q(\x[74][15] ) );
  dp_1 \x_reg[74][14]  ( .ip(n16585), .ck(clk), .q(\x[74][14] ) );
  dp_1 \x_reg[74][13]  ( .ip(n16584), .ck(clk), .q(\x[74][13] ) );
  dp_1 \x_reg[74][12]  ( .ip(n16583), .ck(clk), .q(\x[74][12] ) );
  dp_1 \x_reg[74][11]  ( .ip(n16582), .ck(clk), .q(\x[74][11] ) );
  dp_1 \x_reg[74][10]  ( .ip(n16581), .ck(clk), .q(\x[74][10] ) );
  dp_1 \x_reg[74][9]  ( .ip(n16580), .ck(clk), .q(\x[74][9] ) );
  dp_1 \x_reg[74][8]  ( .ip(n16579), .ck(clk), .q(\x[74][8] ) );
  dp_1 \x_reg[74][7]  ( .ip(n16578), .ck(clk), .q(\x[74][7] ) );
  dp_1 \x_reg[74][6]  ( .ip(n16577), .ck(clk), .q(\x[74][6] ) );
  dp_1 \x_reg[74][5]  ( .ip(n16576), .ck(clk), .q(\x[74][5] ) );
  dp_1 \x_reg[74][4]  ( .ip(n16575), .ck(clk), .q(\x[74][4] ) );
  dp_1 \x_reg[74][3]  ( .ip(n16574), .ck(clk), .q(\x[74][3] ) );
  dp_1 \x_reg[74][2]  ( .ip(n16573), .ck(clk), .q(\x[74][2] ) );
  dp_1 \x_reg[74][1]  ( .ip(n16572), .ck(clk), .q(\x[74][1] ) );
  dp_1 \x_reg[74][0]  ( .ip(n16571), .ck(clk), .q(\x[74][0] ) );
  dp_1 \x_reg[73][15]  ( .ip(n16570), .ck(clk), .q(\x[73][15] ) );
  dp_1 \x_reg[73][14]  ( .ip(n16569), .ck(clk), .q(\x[73][14] ) );
  dp_1 \x_reg[73][13]  ( .ip(n16568), .ck(clk), .q(\x[73][13] ) );
  dp_1 \x_reg[73][12]  ( .ip(n16567), .ck(clk), .q(\x[73][12] ) );
  dp_1 \x_reg[73][11]  ( .ip(n16566), .ck(clk), .q(\x[73][11] ) );
  dp_1 \x_reg[73][10]  ( .ip(n16565), .ck(clk), .q(\x[73][10] ) );
  dp_1 \x_reg[73][9]  ( .ip(n16564), .ck(clk), .q(\x[73][9] ) );
  dp_1 \x_reg[73][8]  ( .ip(n16563), .ck(clk), .q(\x[73][8] ) );
  dp_1 \x_reg[73][7]  ( .ip(n16562), .ck(clk), .q(\x[73][7] ) );
  dp_1 \x_reg[73][6]  ( .ip(n16561), .ck(clk), .q(\x[73][6] ) );
  dp_1 \x_reg[73][5]  ( .ip(n16560), .ck(clk), .q(\x[73][5] ) );
  dp_1 \x_reg[73][4]  ( .ip(n16559), .ck(clk), .q(\x[73][4] ) );
  dp_1 \x_reg[73][3]  ( .ip(n16558), .ck(clk), .q(\x[73][3] ) );
  dp_1 \x_reg[73][2]  ( .ip(n16557), .ck(clk), .q(\x[73][2] ) );
  dp_1 \x_reg[73][1]  ( .ip(n16556), .ck(clk), .q(\x[73][1] ) );
  dp_1 \x_reg[73][0]  ( .ip(n16555), .ck(clk), .q(\x[73][0] ) );
  dp_1 \x_reg[72][15]  ( .ip(n16554), .ck(clk), .q(\x[72][15] ) );
  dp_1 \x_reg[72][14]  ( .ip(n16553), .ck(clk), .q(\x[72][14] ) );
  dp_1 \x_reg[72][13]  ( .ip(n16552), .ck(clk), .q(\x[72][13] ) );
  dp_1 \x_reg[72][12]  ( .ip(n16551), .ck(clk), .q(\x[72][12] ) );
  dp_1 \x_reg[72][11]  ( .ip(n16550), .ck(clk), .q(\x[72][11] ) );
  dp_1 \x_reg[72][10]  ( .ip(n16549), .ck(clk), .q(\x[72][10] ) );
  dp_1 \x_reg[72][9]  ( .ip(n16548), .ck(clk), .q(\x[72][9] ) );
  dp_1 \x_reg[72][8]  ( .ip(n16547), .ck(clk), .q(\x[72][8] ) );
  dp_1 \x_reg[72][7]  ( .ip(n16546), .ck(clk), .q(\x[72][7] ) );
  dp_1 \x_reg[72][6]  ( .ip(n16545), .ck(clk), .q(\x[72][6] ) );
  dp_1 \x_reg[72][5]  ( .ip(n16544), .ck(clk), .q(\x[72][5] ) );
  dp_1 \x_reg[72][4]  ( .ip(n16543), .ck(clk), .q(\x[72][4] ) );
  dp_1 \x_reg[72][3]  ( .ip(n16542), .ck(clk), .q(\x[72][3] ) );
  dp_1 \x_reg[72][2]  ( .ip(n16541), .ck(clk), .q(\x[72][2] ) );
  dp_1 \x_reg[72][1]  ( .ip(n16540), .ck(clk), .q(\x[72][1] ) );
  dp_1 \x_reg[72][0]  ( .ip(n16539), .ck(clk), .q(\x[72][0] ) );
  dp_1 \x_reg[71][15]  ( .ip(n16538), .ck(clk), .q(\x[71][15] ) );
  dp_1 \x_reg[71][14]  ( .ip(n16537), .ck(clk), .q(\x[71][14] ) );
  dp_1 \x_reg[71][13]  ( .ip(n16536), .ck(clk), .q(\x[71][13] ) );
  dp_1 \x_reg[71][12]  ( .ip(n16535), .ck(clk), .q(\x[71][12] ) );
  dp_1 \x_reg[71][11]  ( .ip(n16534), .ck(clk), .q(\x[71][11] ) );
  dp_1 \x_reg[71][10]  ( .ip(n16533), .ck(clk), .q(\x[71][10] ) );
  dp_1 \x_reg[71][9]  ( .ip(n16532), .ck(clk), .q(\x[71][9] ) );
  dp_1 \x_reg[71][8]  ( .ip(n16531), .ck(clk), .q(\x[71][8] ) );
  dp_1 \x_reg[71][7]  ( .ip(n16530), .ck(clk), .q(\x[71][7] ) );
  dp_1 \x_reg[71][6]  ( .ip(n16529), .ck(clk), .q(\x[71][6] ) );
  dp_1 \x_reg[71][5]  ( .ip(n16528), .ck(clk), .q(\x[71][5] ) );
  dp_1 \x_reg[71][4]  ( .ip(n16527), .ck(clk), .q(\x[71][4] ) );
  dp_1 \x_reg[71][3]  ( .ip(n16526), .ck(clk), .q(\x[71][3] ) );
  dp_1 \x_reg[71][2]  ( .ip(n16525), .ck(clk), .q(\x[71][2] ) );
  dp_1 \x_reg[71][1]  ( .ip(n16524), .ck(clk), .q(\x[71][1] ) );
  dp_1 \x_reg[71][0]  ( .ip(n16523), .ck(clk), .q(\x[71][0] ) );
  dp_1 \x_reg[70][15]  ( .ip(n16522), .ck(clk), .q(\x[70][15] ) );
  dp_1 \x_reg[70][14]  ( .ip(n16521), .ck(clk), .q(\x[70][14] ) );
  dp_1 \x_reg[70][13]  ( .ip(n16520), .ck(clk), .q(\x[70][13] ) );
  dp_1 \x_reg[70][12]  ( .ip(n16519), .ck(clk), .q(\x[70][12] ) );
  dp_1 \x_reg[70][11]  ( .ip(n16518), .ck(clk), .q(\x[70][11] ) );
  dp_1 \x_reg[70][10]  ( .ip(n16517), .ck(clk), .q(\x[70][10] ) );
  dp_1 \x_reg[70][9]  ( .ip(n16516), .ck(clk), .q(\x[70][9] ) );
  dp_1 \x_reg[70][8]  ( .ip(n16515), .ck(clk), .q(\x[70][8] ) );
  dp_1 \x_reg[70][7]  ( .ip(n16514), .ck(clk), .q(\x[70][7] ) );
  dp_1 \x_reg[70][6]  ( .ip(n16513), .ck(clk), .q(\x[70][6] ) );
  dp_1 \x_reg[70][5]  ( .ip(n16512), .ck(clk), .q(\x[70][5] ) );
  dp_1 \x_reg[70][4]  ( .ip(n16511), .ck(clk), .q(\x[70][4] ) );
  dp_1 \x_reg[70][3]  ( .ip(n16510), .ck(clk), .q(\x[70][3] ) );
  dp_1 \x_reg[70][2]  ( .ip(n16509), .ck(clk), .q(\x[70][2] ) );
  dp_1 \x_reg[70][1]  ( .ip(n16508), .ck(clk), .q(\x[70][1] ) );
  dp_1 \x_reg[70][0]  ( .ip(n16507), .ck(clk), .q(\x[70][0] ) );
  dp_1 \x_reg[69][15]  ( .ip(n16506), .ck(clk), .q(\x[69][15] ) );
  dp_1 \x_reg[69][14]  ( .ip(n16505), .ck(clk), .q(\x[69][14] ) );
  dp_1 \x_reg[69][13]  ( .ip(n16504), .ck(clk), .q(\x[69][13] ) );
  dp_1 \x_reg[69][12]  ( .ip(n16503), .ck(clk), .q(\x[69][12] ) );
  dp_1 \x_reg[69][11]  ( .ip(n16502), .ck(clk), .q(\x[69][11] ) );
  dp_1 \x_reg[69][10]  ( .ip(n16501), .ck(clk), .q(\x[69][10] ) );
  dp_1 \x_reg[69][9]  ( .ip(n16500), .ck(clk), .q(\x[69][9] ) );
  dp_1 \x_reg[69][8]  ( .ip(n16499), .ck(clk), .q(\x[69][8] ) );
  dp_1 \x_reg[69][7]  ( .ip(n16498), .ck(clk), .q(\x[69][7] ) );
  dp_1 \x_reg[69][6]  ( .ip(n16497), .ck(clk), .q(\x[69][6] ) );
  dp_1 \x_reg[69][5]  ( .ip(n16496), .ck(clk), .q(\x[69][5] ) );
  dp_1 \x_reg[69][4]  ( .ip(n16495), .ck(clk), .q(\x[69][4] ) );
  dp_1 \x_reg[69][3]  ( .ip(n16494), .ck(clk), .q(\x[69][3] ) );
  dp_1 \x_reg[69][2]  ( .ip(n16493), .ck(clk), .q(\x[69][2] ) );
  dp_1 \x_reg[69][1]  ( .ip(n16492), .ck(clk), .q(\x[69][1] ) );
  dp_1 \x_reg[69][0]  ( .ip(n16491), .ck(clk), .q(\x[69][0] ) );
  dp_1 \x_reg[68][15]  ( .ip(n16490), .ck(clk), .q(\x[68][15] ) );
  dp_1 \x_reg[68][14]  ( .ip(n16489), .ck(clk), .q(\x[68][14] ) );
  dp_1 \x_reg[68][13]  ( .ip(n16488), .ck(clk), .q(\x[68][13] ) );
  dp_1 \x_reg[68][12]  ( .ip(n16487), .ck(clk), .q(\x[68][12] ) );
  dp_1 \x_reg[68][11]  ( .ip(n16486), .ck(clk), .q(\x[68][11] ) );
  dp_1 \x_reg[68][10]  ( .ip(n16485), .ck(clk), .q(\x[68][10] ) );
  dp_1 \x_reg[68][9]  ( .ip(n16484), .ck(clk), .q(\x[68][9] ) );
  dp_1 \x_reg[68][8]  ( .ip(n16483), .ck(clk), .q(\x[68][8] ) );
  dp_1 \x_reg[68][7]  ( .ip(n16482), .ck(clk), .q(\x[68][7] ) );
  dp_1 \x_reg[68][6]  ( .ip(n16481), .ck(clk), .q(\x[68][6] ) );
  dp_1 \x_reg[68][5]  ( .ip(n16480), .ck(clk), .q(\x[68][5] ) );
  dp_1 \x_reg[68][4]  ( .ip(n16479), .ck(clk), .q(\x[68][4] ) );
  dp_1 \x_reg[68][3]  ( .ip(n16478), .ck(clk), .q(\x[68][3] ) );
  dp_1 \x_reg[68][2]  ( .ip(n16477), .ck(clk), .q(\x[68][2] ) );
  dp_1 \x_reg[68][1]  ( .ip(n16476), .ck(clk), .q(\x[68][1] ) );
  dp_1 \x_reg[68][0]  ( .ip(n16475), .ck(clk), .q(\x[68][0] ) );
  dp_1 \x_reg[67][15]  ( .ip(n16474), .ck(clk), .q(\x[67][15] ) );
  dp_1 \x_reg[67][14]  ( .ip(n16473), .ck(clk), .q(\x[67][14] ) );
  dp_1 \x_reg[67][13]  ( .ip(n16472), .ck(clk), .q(\x[67][13] ) );
  dp_1 \x_reg[67][12]  ( .ip(n16471), .ck(clk), .q(\x[67][12] ) );
  dp_1 \x_reg[67][11]  ( .ip(n16470), .ck(clk), .q(\x[67][11] ) );
  dp_1 \x_reg[67][10]  ( .ip(n16469), .ck(clk), .q(\x[67][10] ) );
  dp_1 \x_reg[67][9]  ( .ip(n16468), .ck(clk), .q(\x[67][9] ) );
  dp_1 \x_reg[67][8]  ( .ip(n16467), .ck(clk), .q(\x[67][8] ) );
  dp_1 \x_reg[67][7]  ( .ip(n16466), .ck(clk), .q(\x[67][7] ) );
  dp_1 \x_reg[67][6]  ( .ip(n16465), .ck(clk), .q(\x[67][6] ) );
  dp_1 \x_reg[67][5]  ( .ip(n16464), .ck(clk), .q(\x[67][5] ) );
  dp_1 \x_reg[67][4]  ( .ip(n16463), .ck(clk), .q(\x[67][4] ) );
  dp_1 \x_reg[67][3]  ( .ip(n16462), .ck(clk), .q(\x[67][3] ) );
  dp_1 \x_reg[67][2]  ( .ip(n16461), .ck(clk), .q(\x[67][2] ) );
  dp_1 \x_reg[67][1]  ( .ip(n16460), .ck(clk), .q(\x[67][1] ) );
  dp_1 \x_reg[67][0]  ( .ip(n16459), .ck(clk), .q(\x[67][0] ) );
  dp_1 \x_reg[66][15]  ( .ip(n16458), .ck(clk), .q(\x[66][15] ) );
  dp_1 \x_reg[66][14]  ( .ip(n16457), .ck(clk), .q(\x[66][14] ) );
  dp_1 \x_reg[66][13]  ( .ip(n16456), .ck(clk), .q(\x[66][13] ) );
  dp_1 \x_reg[66][12]  ( .ip(n16455), .ck(clk), .q(\x[66][12] ) );
  dp_1 \x_reg[66][11]  ( .ip(n16454), .ck(clk), .q(\x[66][11] ) );
  dp_1 \x_reg[66][10]  ( .ip(n16453), .ck(clk), .q(\x[66][10] ) );
  dp_1 \x_reg[66][9]  ( .ip(n16452), .ck(clk), .q(\x[66][9] ) );
  dp_1 \x_reg[66][8]  ( .ip(n16451), .ck(clk), .q(\x[66][8] ) );
  dp_1 \x_reg[66][7]  ( .ip(n16450), .ck(clk), .q(\x[66][7] ) );
  dp_1 \x_reg[66][6]  ( .ip(n16449), .ck(clk), .q(\x[66][6] ) );
  dp_1 \x_reg[66][5]  ( .ip(n16448), .ck(clk), .q(\x[66][5] ) );
  dp_1 \x_reg[66][4]  ( .ip(n16447), .ck(clk), .q(\x[66][4] ) );
  dp_1 \x_reg[66][3]  ( .ip(n16446), .ck(clk), .q(\x[66][3] ) );
  dp_1 \x_reg[66][2]  ( .ip(n16445), .ck(clk), .q(\x[66][2] ) );
  dp_1 \x_reg[66][1]  ( .ip(n16444), .ck(clk), .q(\x[66][1] ) );
  dp_1 \x_reg[66][0]  ( .ip(n16443), .ck(clk), .q(\x[66][0] ) );
  dp_1 \x_reg[65][15]  ( .ip(n16442), .ck(clk), .q(\x[65][15] ) );
  dp_1 \x_reg[65][14]  ( .ip(n16441), .ck(clk), .q(\x[65][14] ) );
  dp_1 \x_reg[65][13]  ( .ip(n16440), .ck(clk), .q(\x[65][13] ) );
  dp_1 \x_reg[65][12]  ( .ip(n16439), .ck(clk), .q(\x[65][12] ) );
  dp_1 \x_reg[65][11]  ( .ip(n16438), .ck(clk), .q(\x[65][11] ) );
  dp_1 \x_reg[65][10]  ( .ip(n16437), .ck(clk), .q(\x[65][10] ) );
  dp_1 \x_reg[65][9]  ( .ip(n16436), .ck(clk), .q(\x[65][9] ) );
  dp_1 \x_reg[65][8]  ( .ip(n16435), .ck(clk), .q(\x[65][8] ) );
  dp_1 \x_reg[65][7]  ( .ip(n16434), .ck(clk), .q(\x[65][7] ) );
  dp_1 \x_reg[65][6]  ( .ip(n16433), .ck(clk), .q(\x[65][6] ) );
  dp_1 \x_reg[65][5]  ( .ip(n16432), .ck(clk), .q(\x[65][5] ) );
  dp_1 \x_reg[65][4]  ( .ip(n16431), .ck(clk), .q(\x[65][4] ) );
  dp_1 \x_reg[65][3]  ( .ip(n16430), .ck(clk), .q(\x[65][3] ) );
  dp_1 \x_reg[65][2]  ( .ip(n16429), .ck(clk), .q(\x[65][2] ) );
  dp_1 \x_reg[65][1]  ( .ip(n16428), .ck(clk), .q(\x[65][1] ) );
  dp_1 \x_reg[65][0]  ( .ip(n16427), .ck(clk), .q(\x[65][0] ) );
  dp_1 \x_reg[64][15]  ( .ip(n16426), .ck(clk), .q(\x[64][15] ) );
  dp_1 \x_reg[64][14]  ( .ip(n16425), .ck(clk), .q(\x[64][14] ) );
  dp_1 \x_reg[64][13]  ( .ip(n16424), .ck(clk), .q(\x[64][13] ) );
  dp_1 \x_reg[64][12]  ( .ip(n16423), .ck(clk), .q(\x[64][12] ) );
  dp_1 \x_reg[64][11]  ( .ip(n16422), .ck(clk), .q(\x[64][11] ) );
  dp_1 \x_reg[64][10]  ( .ip(n16421), .ck(clk), .q(\x[64][10] ) );
  dp_1 \x_reg[64][9]  ( .ip(n16420), .ck(clk), .q(\x[64][9] ) );
  dp_1 \x_reg[64][8]  ( .ip(n16419), .ck(clk), .q(\x[64][8] ) );
  dp_1 \x_reg[64][7]  ( .ip(n16418), .ck(clk), .q(\x[64][7] ) );
  dp_1 \x_reg[64][6]  ( .ip(n16417), .ck(clk), .q(\x[64][6] ) );
  dp_1 \x_reg[64][5]  ( .ip(n16416), .ck(clk), .q(\x[64][5] ) );
  dp_1 \x_reg[64][4]  ( .ip(n16415), .ck(clk), .q(\x[64][4] ) );
  dp_1 \x_reg[64][3]  ( .ip(n16414), .ck(clk), .q(\x[64][3] ) );
  dp_1 \x_reg[64][2]  ( .ip(n16413), .ck(clk), .q(\x[64][2] ) );
  dp_1 \x_reg[64][1]  ( .ip(n16412), .ck(clk), .q(\x[64][1] ) );
  dp_1 \x_reg[64][0]  ( .ip(n16411), .ck(clk), .q(\x[64][0] ) );
  dp_1 \x_reg[63][15]  ( .ip(n16410), .ck(clk), .q(\x[63][15] ) );
  dp_1 \x_reg[63][14]  ( .ip(n16409), .ck(clk), .q(\x[63][14] ) );
  dp_1 \x_reg[63][13]  ( .ip(n16408), .ck(clk), .q(\x[63][13] ) );
  dp_1 \x_reg[63][12]  ( .ip(n16407), .ck(clk), .q(\x[63][12] ) );
  dp_1 \x_reg[63][11]  ( .ip(n16406), .ck(clk), .q(\x[63][11] ) );
  dp_1 \x_reg[63][10]  ( .ip(n16405), .ck(clk), .q(\x[63][10] ) );
  dp_1 \x_reg[63][9]  ( .ip(n16404), .ck(clk), .q(\x[63][9] ) );
  dp_1 \x_reg[63][8]  ( .ip(n16403), .ck(clk), .q(\x[63][8] ) );
  dp_1 \x_reg[63][7]  ( .ip(n16402), .ck(clk), .q(\x[63][7] ) );
  dp_1 \x_reg[63][6]  ( .ip(n16401), .ck(clk), .q(\x[63][6] ) );
  dp_1 \x_reg[63][5]  ( .ip(n16400), .ck(clk), .q(\x[63][5] ) );
  dp_1 \x_reg[63][4]  ( .ip(n16399), .ck(clk), .q(\x[63][4] ) );
  dp_1 \x_reg[63][3]  ( .ip(n16398), .ck(clk), .q(\x[63][3] ) );
  dp_1 \x_reg[63][2]  ( .ip(n16397), .ck(clk), .q(\x[63][2] ) );
  dp_1 \x_reg[63][1]  ( .ip(n16396), .ck(clk), .q(\x[63][1] ) );
  dp_1 \x_reg[63][0]  ( .ip(n16395), .ck(clk), .q(\x[63][0] ) );
  dp_1 \x_reg[62][15]  ( .ip(n16394), .ck(clk), .q(\x[62][15] ) );
  dp_1 \x_reg[62][14]  ( .ip(n16393), .ck(clk), .q(\x[62][14] ) );
  dp_1 \x_reg[62][13]  ( .ip(n16392), .ck(clk), .q(\x[62][13] ) );
  dp_1 \x_reg[62][12]  ( .ip(n16391), .ck(clk), .q(\x[62][12] ) );
  dp_1 \x_reg[62][11]  ( .ip(n16390), .ck(clk), .q(\x[62][11] ) );
  dp_1 \x_reg[62][10]  ( .ip(n16389), .ck(clk), .q(\x[62][10] ) );
  dp_1 \x_reg[62][9]  ( .ip(n16388), .ck(clk), .q(\x[62][9] ) );
  dp_1 \x_reg[62][8]  ( .ip(n16387), .ck(clk), .q(\x[62][8] ) );
  dp_1 \x_reg[62][7]  ( .ip(n16386), .ck(clk), .q(\x[62][7] ) );
  dp_1 \x_reg[62][6]  ( .ip(n16385), .ck(clk), .q(\x[62][6] ) );
  dp_1 \x_reg[62][5]  ( .ip(n16384), .ck(clk), .q(\x[62][5] ) );
  dp_1 \x_reg[62][4]  ( .ip(n16383), .ck(clk), .q(\x[62][4] ) );
  dp_1 \x_reg[62][3]  ( .ip(n16382), .ck(clk), .q(\x[62][3] ) );
  dp_1 \x_reg[62][2]  ( .ip(n16381), .ck(clk), .q(\x[62][2] ) );
  dp_1 \x_reg[62][1]  ( .ip(n16380), .ck(clk), .q(\x[62][1] ) );
  dp_1 \x_reg[62][0]  ( .ip(n16379), .ck(clk), .q(\x[62][0] ) );
  dp_1 \x_reg[61][15]  ( .ip(n16378), .ck(clk), .q(\x[61][15] ) );
  dp_1 \x_reg[61][14]  ( .ip(n16377), .ck(clk), .q(\x[61][14] ) );
  dp_1 \x_reg[61][13]  ( .ip(n16376), .ck(clk), .q(\x[61][13] ) );
  dp_1 \x_reg[61][12]  ( .ip(n16375), .ck(clk), .q(\x[61][12] ) );
  dp_1 \x_reg[61][11]  ( .ip(n16374), .ck(clk), .q(\x[61][11] ) );
  dp_1 \x_reg[61][10]  ( .ip(n16373), .ck(clk), .q(\x[61][10] ) );
  dp_1 \x_reg[61][9]  ( .ip(n16372), .ck(clk), .q(\x[61][9] ) );
  dp_1 \x_reg[61][8]  ( .ip(n16371), .ck(clk), .q(\x[61][8] ) );
  dp_1 \x_reg[61][7]  ( .ip(n16370), .ck(clk), .q(\x[61][7] ) );
  dp_1 \x_reg[61][6]  ( .ip(n16369), .ck(clk), .q(\x[61][6] ) );
  dp_1 \x_reg[61][5]  ( .ip(n16368), .ck(clk), .q(\x[61][5] ) );
  dp_1 \x_reg[61][4]  ( .ip(n16367), .ck(clk), .q(\x[61][4] ) );
  dp_1 \x_reg[61][3]  ( .ip(n16366), .ck(clk), .q(\x[61][3] ) );
  dp_1 \x_reg[61][2]  ( .ip(n16365), .ck(clk), .q(\x[61][2] ) );
  dp_1 \x_reg[61][1]  ( .ip(n16364), .ck(clk), .q(\x[61][1] ) );
  dp_1 \x_reg[61][0]  ( .ip(n16363), .ck(clk), .q(\x[61][0] ) );
  dp_1 \x_reg[60][15]  ( .ip(n16362), .ck(clk), .q(\x[60][15] ) );
  dp_1 \x_reg[60][14]  ( .ip(n16361), .ck(clk), .q(\x[60][14] ) );
  dp_1 \x_reg[60][13]  ( .ip(n16360), .ck(clk), .q(\x[60][13] ) );
  dp_1 \x_reg[60][12]  ( .ip(n16359), .ck(clk), .q(\x[60][12] ) );
  dp_1 \x_reg[60][11]  ( .ip(n16358), .ck(clk), .q(\x[60][11] ) );
  dp_1 \x_reg[60][10]  ( .ip(n16357), .ck(clk), .q(\x[60][10] ) );
  dp_1 \x_reg[60][9]  ( .ip(n16356), .ck(clk), .q(\x[60][9] ) );
  dp_1 \x_reg[60][8]  ( .ip(n16355), .ck(clk), .q(\x[60][8] ) );
  dp_1 \x_reg[60][7]  ( .ip(n16354), .ck(clk), .q(\x[60][7] ) );
  dp_1 \x_reg[60][6]  ( .ip(n16353), .ck(clk), .q(\x[60][6] ) );
  dp_1 \x_reg[60][5]  ( .ip(n16352), .ck(clk), .q(\x[60][5] ) );
  dp_1 \x_reg[60][4]  ( .ip(n16351), .ck(clk), .q(\x[60][4] ) );
  dp_1 \x_reg[60][3]  ( .ip(n16350), .ck(clk), .q(\x[60][3] ) );
  dp_1 \x_reg[60][2]  ( .ip(n16349), .ck(clk), .q(\x[60][2] ) );
  dp_1 \x_reg[60][1]  ( .ip(n16348), .ck(clk), .q(\x[60][1] ) );
  dp_1 \x_reg[60][0]  ( .ip(n16347), .ck(clk), .q(\x[60][0] ) );
  dp_1 \x_reg[59][15]  ( .ip(n16346), .ck(clk), .q(\x[59][15] ) );
  dp_1 \x_reg[59][14]  ( .ip(n16345), .ck(clk), .q(\x[59][14] ) );
  dp_1 \x_reg[59][13]  ( .ip(n16344), .ck(clk), .q(\x[59][13] ) );
  dp_1 \x_reg[59][12]  ( .ip(n16343), .ck(clk), .q(\x[59][12] ) );
  dp_1 \x_reg[59][11]  ( .ip(n16342), .ck(clk), .q(\x[59][11] ) );
  dp_1 \x_reg[59][10]  ( .ip(n16341), .ck(clk), .q(\x[59][10] ) );
  dp_1 \x_reg[59][9]  ( .ip(n16340), .ck(clk), .q(\x[59][9] ) );
  dp_1 \x_reg[59][8]  ( .ip(n16339), .ck(clk), .q(\x[59][8] ) );
  dp_1 \x_reg[59][7]  ( .ip(n16338), .ck(clk), .q(\x[59][7] ) );
  dp_1 \x_reg[59][6]  ( .ip(n16337), .ck(clk), .q(\x[59][6] ) );
  dp_1 \x_reg[59][5]  ( .ip(n16336), .ck(clk), .q(\x[59][5] ) );
  dp_1 \x_reg[59][4]  ( .ip(n16335), .ck(clk), .q(\x[59][4] ) );
  dp_1 \x_reg[59][3]  ( .ip(n16334), .ck(clk), .q(\x[59][3] ) );
  dp_1 \x_reg[59][2]  ( .ip(n16333), .ck(clk), .q(\x[59][2] ) );
  dp_1 \x_reg[59][1]  ( .ip(n16332), .ck(clk), .q(\x[59][1] ) );
  dp_1 \x_reg[59][0]  ( .ip(n16331), .ck(clk), .q(\x[59][0] ) );
  dp_1 \x_reg[58][15]  ( .ip(n16330), .ck(clk), .q(\x[58][15] ) );
  dp_1 \x_reg[58][14]  ( .ip(n16329), .ck(clk), .q(\x[58][14] ) );
  dp_1 \x_reg[58][13]  ( .ip(n16328), .ck(clk), .q(\x[58][13] ) );
  dp_1 \x_reg[58][12]  ( .ip(n16327), .ck(clk), .q(\x[58][12] ) );
  dp_1 \x_reg[58][11]  ( .ip(n16326), .ck(clk), .q(\x[58][11] ) );
  dp_1 \x_reg[58][10]  ( .ip(n16325), .ck(clk), .q(\x[58][10] ) );
  dp_1 \x_reg[58][9]  ( .ip(n16324), .ck(clk), .q(\x[58][9] ) );
  dp_1 \x_reg[58][8]  ( .ip(n16323), .ck(clk), .q(\x[58][8] ) );
  dp_1 \x_reg[58][7]  ( .ip(n16322), .ck(clk), .q(\x[58][7] ) );
  dp_1 \x_reg[58][6]  ( .ip(n16321), .ck(clk), .q(\x[58][6] ) );
  dp_1 \x_reg[58][5]  ( .ip(n16320), .ck(clk), .q(\x[58][5] ) );
  dp_1 \x_reg[58][4]  ( .ip(n16319), .ck(clk), .q(\x[58][4] ) );
  dp_1 \x_reg[58][3]  ( .ip(n16318), .ck(clk), .q(\x[58][3] ) );
  dp_1 \x_reg[58][2]  ( .ip(n16317), .ck(clk), .q(\x[58][2] ) );
  dp_1 \x_reg[58][1]  ( .ip(n16316), .ck(clk), .q(\x[58][1] ) );
  dp_1 \x_reg[58][0]  ( .ip(n16315), .ck(clk), .q(\x[58][0] ) );
  dp_1 \x_reg[57][15]  ( .ip(n16314), .ck(clk), .q(\x[57][15] ) );
  dp_1 \x_reg[57][14]  ( .ip(n16313), .ck(clk), .q(\x[57][14] ) );
  dp_1 \x_reg[57][13]  ( .ip(n16312), .ck(clk), .q(\x[57][13] ) );
  dp_1 \x_reg[57][12]  ( .ip(n16311), .ck(clk), .q(\x[57][12] ) );
  dp_1 \x_reg[57][11]  ( .ip(n16310), .ck(clk), .q(\x[57][11] ) );
  dp_1 \x_reg[57][10]  ( .ip(n16309), .ck(clk), .q(\x[57][10] ) );
  dp_1 \x_reg[57][9]  ( .ip(n16308), .ck(clk), .q(\x[57][9] ) );
  dp_1 \x_reg[57][8]  ( .ip(n16307), .ck(clk), .q(\x[57][8] ) );
  dp_1 \x_reg[57][7]  ( .ip(n16306), .ck(clk), .q(\x[57][7] ) );
  dp_1 \x_reg[57][6]  ( .ip(n16305), .ck(clk), .q(\x[57][6] ) );
  dp_1 \x_reg[57][5]  ( .ip(n16304), .ck(clk), .q(\x[57][5] ) );
  dp_1 \x_reg[57][4]  ( .ip(n16303), .ck(clk), .q(\x[57][4] ) );
  dp_1 \x_reg[57][3]  ( .ip(n16302), .ck(clk), .q(\x[57][3] ) );
  dp_1 \x_reg[57][2]  ( .ip(n16301), .ck(clk), .q(\x[57][2] ) );
  dp_1 \x_reg[57][1]  ( .ip(n16300), .ck(clk), .q(\x[57][1] ) );
  dp_1 \x_reg[57][0]  ( .ip(n16299), .ck(clk), .q(\x[57][0] ) );
  dp_1 \x_reg[56][15]  ( .ip(n16298), .ck(clk), .q(\x[56][15] ) );
  dp_1 \x_reg[56][14]  ( .ip(n16297), .ck(clk), .q(\x[56][14] ) );
  dp_1 \x_reg[56][13]  ( .ip(n16296), .ck(clk), .q(\x[56][13] ) );
  dp_1 \x_reg[56][12]  ( .ip(n16295), .ck(clk), .q(\x[56][12] ) );
  dp_1 \x_reg[56][11]  ( .ip(n16294), .ck(clk), .q(\x[56][11] ) );
  dp_1 \x_reg[56][10]  ( .ip(n16293), .ck(clk), .q(\x[56][10] ) );
  dp_1 \x_reg[56][9]  ( .ip(n16292), .ck(clk), .q(\x[56][9] ) );
  dp_1 \x_reg[56][8]  ( .ip(n16291), .ck(clk), .q(\x[56][8] ) );
  dp_1 \x_reg[56][7]  ( .ip(n16290), .ck(clk), .q(\x[56][7] ) );
  dp_1 \x_reg[56][6]  ( .ip(n16289), .ck(clk), .q(\x[56][6] ) );
  dp_1 \x_reg[56][5]  ( .ip(n16288), .ck(clk), .q(\x[56][5] ) );
  dp_1 \x_reg[56][4]  ( .ip(n16287), .ck(clk), .q(\x[56][4] ) );
  dp_1 \x_reg[56][3]  ( .ip(n16286), .ck(clk), .q(\x[56][3] ) );
  dp_1 \x_reg[56][2]  ( .ip(n16285), .ck(clk), .q(\x[56][2] ) );
  dp_1 \x_reg[56][1]  ( .ip(n16284), .ck(clk), .q(\x[56][1] ) );
  dp_1 \x_reg[56][0]  ( .ip(n16283), .ck(clk), .q(\x[56][0] ) );
  dp_1 \x_reg[55][15]  ( .ip(n16282), .ck(clk), .q(\x[55][15] ) );
  dp_1 \x_reg[55][14]  ( .ip(n16281), .ck(clk), .q(\x[55][14] ) );
  dp_1 \x_reg[55][13]  ( .ip(n16280), .ck(clk), .q(\x[55][13] ) );
  dp_1 \x_reg[55][12]  ( .ip(n16279), .ck(clk), .q(\x[55][12] ) );
  dp_1 \x_reg[55][11]  ( .ip(n16278), .ck(clk), .q(\x[55][11] ) );
  dp_1 \x_reg[55][10]  ( .ip(n16277), .ck(clk), .q(\x[55][10] ) );
  dp_1 \x_reg[55][9]  ( .ip(n16276), .ck(clk), .q(\x[55][9] ) );
  dp_1 \x_reg[55][8]  ( .ip(n16275), .ck(clk), .q(\x[55][8] ) );
  dp_1 \x_reg[55][7]  ( .ip(n16274), .ck(clk), .q(\x[55][7] ) );
  dp_1 \x_reg[55][6]  ( .ip(n16273), .ck(clk), .q(\x[55][6] ) );
  dp_1 \x_reg[55][5]  ( .ip(n16272), .ck(clk), .q(\x[55][5] ) );
  dp_1 \x_reg[55][4]  ( .ip(n16271), .ck(clk), .q(\x[55][4] ) );
  dp_1 \x_reg[55][3]  ( .ip(n16270), .ck(clk), .q(\x[55][3] ) );
  dp_1 \x_reg[55][2]  ( .ip(n16269), .ck(clk), .q(\x[55][2] ) );
  dp_1 \x_reg[55][1]  ( .ip(n16268), .ck(clk), .q(\x[55][1] ) );
  dp_1 \x_reg[55][0]  ( .ip(n16267), .ck(clk), .q(\x[55][0] ) );
  dp_1 \x_reg[54][15]  ( .ip(n16266), .ck(clk), .q(\x[54][15] ) );
  dp_1 \x_reg[54][14]  ( .ip(n16265), .ck(clk), .q(\x[54][14] ) );
  dp_1 \x_reg[54][13]  ( .ip(n16264), .ck(clk), .q(\x[54][13] ) );
  dp_1 \x_reg[54][12]  ( .ip(n16263), .ck(clk), .q(\x[54][12] ) );
  dp_1 \x_reg[54][11]  ( .ip(n16262), .ck(clk), .q(\x[54][11] ) );
  dp_1 \x_reg[54][10]  ( .ip(n16261), .ck(clk), .q(\x[54][10] ) );
  dp_1 \x_reg[54][9]  ( .ip(n16260), .ck(clk), .q(\x[54][9] ) );
  dp_1 \x_reg[54][8]  ( .ip(n16259), .ck(clk), .q(\x[54][8] ) );
  dp_1 \x_reg[54][7]  ( .ip(n16258), .ck(clk), .q(\x[54][7] ) );
  dp_1 \x_reg[54][6]  ( .ip(n16257), .ck(clk), .q(\x[54][6] ) );
  dp_1 \x_reg[54][5]  ( .ip(n16256), .ck(clk), .q(\x[54][5] ) );
  dp_1 \x_reg[54][4]  ( .ip(n16255), .ck(clk), .q(\x[54][4] ) );
  dp_1 \x_reg[54][3]  ( .ip(n16254), .ck(clk), .q(\x[54][3] ) );
  dp_1 \x_reg[54][2]  ( .ip(n16253), .ck(clk), .q(\x[54][2] ) );
  dp_1 \x_reg[54][1]  ( .ip(n16252), .ck(clk), .q(\x[54][1] ) );
  dp_1 \x_reg[54][0]  ( .ip(n16251), .ck(clk), .q(\x[54][0] ) );
  dp_1 \x_reg[53][15]  ( .ip(n16250), .ck(clk), .q(\x[53][15] ) );
  dp_1 \x_reg[53][14]  ( .ip(n16249), .ck(clk), .q(\x[53][14] ) );
  dp_1 \x_reg[53][13]  ( .ip(n16248), .ck(clk), .q(\x[53][13] ) );
  dp_1 \x_reg[53][12]  ( .ip(n16247), .ck(clk), .q(\x[53][12] ) );
  dp_1 \x_reg[53][11]  ( .ip(n16246), .ck(clk), .q(\x[53][11] ) );
  dp_1 \x_reg[53][10]  ( .ip(n16245), .ck(clk), .q(\x[53][10] ) );
  dp_1 \x_reg[53][9]  ( .ip(n16244), .ck(clk), .q(\x[53][9] ) );
  dp_1 \x_reg[53][8]  ( .ip(n16243), .ck(clk), .q(\x[53][8] ) );
  dp_1 \x_reg[53][7]  ( .ip(n16242), .ck(clk), .q(\x[53][7] ) );
  dp_1 \x_reg[53][6]  ( .ip(n16241), .ck(clk), .q(\x[53][6] ) );
  dp_1 \x_reg[53][5]  ( .ip(n16240), .ck(clk), .q(\x[53][5] ) );
  dp_1 \x_reg[53][4]  ( .ip(n16239), .ck(clk), .q(\x[53][4] ) );
  dp_1 \x_reg[53][3]  ( .ip(n16238), .ck(clk), .q(\x[53][3] ) );
  dp_1 \x_reg[53][2]  ( .ip(n16237), .ck(clk), .q(\x[53][2] ) );
  dp_1 \x_reg[53][1]  ( .ip(n16236), .ck(clk), .q(\x[53][1] ) );
  dp_1 \x_reg[53][0]  ( .ip(n16235), .ck(clk), .q(\x[53][0] ) );
  dp_1 \x_reg[52][15]  ( .ip(n16234), .ck(clk), .q(\x[52][15] ) );
  dp_1 \x_reg[52][14]  ( .ip(n16233), .ck(clk), .q(\x[52][14] ) );
  dp_1 \x_reg[52][13]  ( .ip(n16232), .ck(clk), .q(\x[52][13] ) );
  dp_1 \x_reg[52][12]  ( .ip(n16231), .ck(clk), .q(\x[52][12] ) );
  dp_1 \x_reg[52][11]  ( .ip(n16230), .ck(clk), .q(\x[52][11] ) );
  dp_1 \x_reg[52][10]  ( .ip(n16229), .ck(clk), .q(\x[52][10] ) );
  dp_1 \x_reg[52][9]  ( .ip(n16228), .ck(clk), .q(\x[52][9] ) );
  dp_1 \x_reg[52][8]  ( .ip(n16227), .ck(clk), .q(\x[52][8] ) );
  dp_1 \x_reg[52][7]  ( .ip(n16226), .ck(clk), .q(\x[52][7] ) );
  dp_1 \x_reg[52][6]  ( .ip(n16225), .ck(clk), .q(\x[52][6] ) );
  dp_1 \x_reg[52][5]  ( .ip(n16224), .ck(clk), .q(\x[52][5] ) );
  dp_1 \x_reg[52][4]  ( .ip(n16223), .ck(clk), .q(\x[52][4] ) );
  dp_1 \x_reg[52][3]  ( .ip(n16222), .ck(clk), .q(\x[52][3] ) );
  dp_1 \x_reg[52][2]  ( .ip(n16221), .ck(clk), .q(\x[52][2] ) );
  dp_1 \x_reg[52][1]  ( .ip(n16220), .ck(clk), .q(\x[52][1] ) );
  dp_1 \x_reg[52][0]  ( .ip(n16219), .ck(clk), .q(\x[52][0] ) );
  dp_1 \x_reg[51][15]  ( .ip(n16218), .ck(clk), .q(\x[51][15] ) );
  dp_1 \x_reg[51][14]  ( .ip(n16217), .ck(clk), .q(\x[51][14] ) );
  dp_1 \x_reg[51][13]  ( .ip(n16216), .ck(clk), .q(\x[51][13] ) );
  dp_1 \x_reg[51][12]  ( .ip(n16215), .ck(clk), .q(\x[51][12] ) );
  dp_1 \x_reg[51][11]  ( .ip(n16214), .ck(clk), .q(\x[51][11] ) );
  dp_1 \x_reg[51][10]  ( .ip(n16213), .ck(clk), .q(\x[51][10] ) );
  dp_1 \x_reg[51][9]  ( .ip(n16212), .ck(clk), .q(\x[51][9] ) );
  dp_1 \x_reg[51][8]  ( .ip(n16211), .ck(clk), .q(\x[51][8] ) );
  dp_1 \x_reg[51][7]  ( .ip(n16210), .ck(clk), .q(\x[51][7] ) );
  dp_1 \x_reg[51][6]  ( .ip(n16209), .ck(clk), .q(\x[51][6] ) );
  dp_1 \x_reg[51][5]  ( .ip(n16208), .ck(clk), .q(\x[51][5] ) );
  dp_1 \x_reg[51][4]  ( .ip(n16207), .ck(clk), .q(\x[51][4] ) );
  dp_1 \x_reg[51][3]  ( .ip(n16206), .ck(clk), .q(\x[51][3] ) );
  dp_1 \x_reg[51][2]  ( .ip(n16205), .ck(clk), .q(\x[51][2] ) );
  dp_1 \x_reg[51][1]  ( .ip(n16204), .ck(clk), .q(\x[51][1] ) );
  dp_1 \x_reg[51][0]  ( .ip(n16203), .ck(clk), .q(\x[51][0] ) );
  dp_1 \x_reg[50][15]  ( .ip(n16202), .ck(clk), .q(\x[50][15] ) );
  dp_1 \x_reg[50][14]  ( .ip(n16201), .ck(clk), .q(\x[50][14] ) );
  dp_1 \x_reg[50][13]  ( .ip(n16200), .ck(clk), .q(\x[50][13] ) );
  dp_1 \x_reg[50][12]  ( .ip(n16199), .ck(clk), .q(\x[50][12] ) );
  dp_1 \x_reg[50][11]  ( .ip(n16198), .ck(clk), .q(\x[50][11] ) );
  dp_1 \x_reg[50][10]  ( .ip(n16197), .ck(clk), .q(\x[50][10] ) );
  dp_1 \x_reg[50][9]  ( .ip(n16196), .ck(clk), .q(\x[50][9] ) );
  dp_1 \x_reg[50][8]  ( .ip(n16195), .ck(clk), .q(\x[50][8] ) );
  dp_1 \x_reg[50][7]  ( .ip(n16194), .ck(clk), .q(\x[50][7] ) );
  dp_1 \x_reg[50][6]  ( .ip(n16193), .ck(clk), .q(\x[50][6] ) );
  dp_1 \x_reg[50][5]  ( .ip(n16192), .ck(clk), .q(\x[50][5] ) );
  dp_1 \x_reg[50][4]  ( .ip(n16191), .ck(clk), .q(\x[50][4] ) );
  dp_1 \x_reg[50][3]  ( .ip(n16190), .ck(clk), .q(\x[50][3] ) );
  dp_1 \x_reg[50][2]  ( .ip(n16189), .ck(clk), .q(\x[50][2] ) );
  dp_1 \x_reg[50][1]  ( .ip(n16188), .ck(clk), .q(\x[50][1] ) );
  dp_1 \x_reg[50][0]  ( .ip(n16187), .ck(clk), .q(\x[50][0] ) );
  dp_1 \x_reg[49][15]  ( .ip(n16186), .ck(clk), .q(\x[49][15] ) );
  dp_1 \x_reg[49][14]  ( .ip(n16185), .ck(clk), .q(\x[49][14] ) );
  dp_1 \x_reg[49][13]  ( .ip(n16184), .ck(clk), .q(\x[49][13] ) );
  dp_1 \x_reg[49][12]  ( .ip(n16183), .ck(clk), .q(\x[49][12] ) );
  dp_1 \x_reg[49][11]  ( .ip(n16182), .ck(clk), .q(\x[49][11] ) );
  dp_1 \x_reg[49][10]  ( .ip(n16181), .ck(clk), .q(\x[49][10] ) );
  dp_1 \x_reg[49][9]  ( .ip(n16180), .ck(clk), .q(\x[49][9] ) );
  dp_1 \x_reg[49][8]  ( .ip(n16179), .ck(clk), .q(\x[49][8] ) );
  dp_1 \x_reg[49][7]  ( .ip(n16178), .ck(clk), .q(\x[49][7] ) );
  dp_1 \x_reg[49][6]  ( .ip(n16177), .ck(clk), .q(\x[49][6] ) );
  dp_1 \x_reg[49][5]  ( .ip(n16176), .ck(clk), .q(\x[49][5] ) );
  dp_1 \x_reg[49][4]  ( .ip(n16175), .ck(clk), .q(\x[49][4] ) );
  dp_1 \x_reg[49][3]  ( .ip(n16174), .ck(clk), .q(\x[49][3] ) );
  dp_1 \x_reg[49][2]  ( .ip(n16173), .ck(clk), .q(\x[49][2] ) );
  dp_1 \x_reg[49][1]  ( .ip(n16172), .ck(clk), .q(\x[49][1] ) );
  dp_1 \x_reg[49][0]  ( .ip(n16171), .ck(clk), .q(\x[49][0] ) );
  dp_1 \x_reg[48][15]  ( .ip(n16170), .ck(clk), .q(\x[48][15] ) );
  dp_1 \x_reg[48][14]  ( .ip(n16169), .ck(clk), .q(\x[48][14] ) );
  dp_1 \x_reg[48][13]  ( .ip(n16168), .ck(clk), .q(\x[48][13] ) );
  dp_1 \x_reg[48][12]  ( .ip(n16167), .ck(clk), .q(\x[48][12] ) );
  dp_1 \x_reg[48][11]  ( .ip(n16166), .ck(clk), .q(\x[48][11] ) );
  dp_1 \x_reg[48][10]  ( .ip(n16165), .ck(clk), .q(\x[48][10] ) );
  dp_1 \x_reg[48][9]  ( .ip(n16164), .ck(clk), .q(\x[48][9] ) );
  dp_1 \x_reg[48][8]  ( .ip(n16163), .ck(clk), .q(\x[48][8] ) );
  dp_1 \x_reg[48][7]  ( .ip(n16162), .ck(clk), .q(\x[48][7] ) );
  dp_1 \x_reg[48][6]  ( .ip(n16161), .ck(clk), .q(\x[48][6] ) );
  dp_1 \x_reg[48][5]  ( .ip(n16160), .ck(clk), .q(\x[48][5] ) );
  dp_1 \x_reg[48][4]  ( .ip(n16159), .ck(clk), .q(\x[48][4] ) );
  dp_1 \x_reg[48][3]  ( .ip(n16158), .ck(clk), .q(\x[48][3] ) );
  dp_1 \x_reg[48][2]  ( .ip(n16157), .ck(clk), .q(\x[48][2] ) );
  dp_1 \x_reg[48][1]  ( .ip(n16156), .ck(clk), .q(\x[48][1] ) );
  dp_1 \x_reg[48][0]  ( .ip(n16155), .ck(clk), .q(\x[48][0] ) );
  dp_1 \x_reg[47][15]  ( .ip(n16154), .ck(clk), .q(\x[47][15] ) );
  dp_1 \x_reg[47][14]  ( .ip(n16153), .ck(clk), .q(\x[47][14] ) );
  dp_1 \x_reg[47][13]  ( .ip(n16152), .ck(clk), .q(\x[47][13] ) );
  dp_1 \x_reg[47][12]  ( .ip(n16151), .ck(clk), .q(\x[47][12] ) );
  dp_1 \x_reg[47][11]  ( .ip(n16150), .ck(clk), .q(\x[47][11] ) );
  dp_1 \x_reg[47][10]  ( .ip(n16149), .ck(clk), .q(\x[47][10] ) );
  dp_1 \x_reg[47][9]  ( .ip(n16148), .ck(clk), .q(\x[47][9] ) );
  dp_1 \x_reg[47][8]  ( .ip(n16147), .ck(clk), .q(\x[47][8] ) );
  dp_1 \x_reg[47][7]  ( .ip(n16146), .ck(clk), .q(\x[47][7] ) );
  dp_1 \x_reg[47][6]  ( .ip(n16145), .ck(clk), .q(\x[47][6] ) );
  dp_1 \x_reg[47][5]  ( .ip(n16144), .ck(clk), .q(\x[47][5] ) );
  dp_1 \x_reg[47][4]  ( .ip(n16143), .ck(clk), .q(\x[47][4] ) );
  dp_1 \x_reg[47][3]  ( .ip(n16142), .ck(clk), .q(\x[47][3] ) );
  dp_1 \x_reg[47][2]  ( .ip(n16141), .ck(clk), .q(\x[47][2] ) );
  dp_1 \x_reg[47][1]  ( .ip(n16140), .ck(clk), .q(\x[47][1] ) );
  dp_1 \x_reg[47][0]  ( .ip(n16139), .ck(clk), .q(\x[47][0] ) );
  dp_1 \x_reg[46][15]  ( .ip(n16138), .ck(clk), .q(\x[46][15] ) );
  dp_1 \x_reg[46][14]  ( .ip(n16137), .ck(clk), .q(\x[46][14] ) );
  dp_1 \x_reg[46][13]  ( .ip(n16136), .ck(clk), .q(\x[46][13] ) );
  dp_1 \x_reg[46][12]  ( .ip(n16135), .ck(clk), .q(\x[46][12] ) );
  dp_1 \x_reg[46][11]  ( .ip(n16134), .ck(clk), .q(\x[46][11] ) );
  dp_1 \x_reg[46][10]  ( .ip(n16133), .ck(clk), .q(\x[46][10] ) );
  dp_1 \x_reg[46][9]  ( .ip(n16132), .ck(clk), .q(\x[46][9] ) );
  dp_1 \x_reg[46][8]  ( .ip(n16131), .ck(clk), .q(\x[46][8] ) );
  dp_1 \x_reg[46][7]  ( .ip(n16130), .ck(clk), .q(\x[46][7] ) );
  dp_1 \x_reg[46][6]  ( .ip(n16129), .ck(clk), .q(\x[46][6] ) );
  dp_1 \x_reg[46][5]  ( .ip(n16128), .ck(clk), .q(\x[46][5] ) );
  dp_1 \x_reg[46][4]  ( .ip(n16127), .ck(clk), .q(\x[46][4] ) );
  dp_1 \x_reg[46][3]  ( .ip(n16126), .ck(clk), .q(\x[46][3] ) );
  dp_1 \x_reg[46][2]  ( .ip(n16125), .ck(clk), .q(\x[46][2] ) );
  dp_1 \x_reg[46][1]  ( .ip(n16124), .ck(clk), .q(\x[46][1] ) );
  dp_1 \x_reg[46][0]  ( .ip(n16123), .ck(clk), .q(\x[46][0] ) );
  dp_1 \x_reg[45][15]  ( .ip(n16122), .ck(clk), .q(\x[45][15] ) );
  dp_1 \x_reg[45][14]  ( .ip(n16121), .ck(clk), .q(\x[45][14] ) );
  dp_1 \x_reg[45][13]  ( .ip(n16120), .ck(clk), .q(\x[45][13] ) );
  dp_1 \x_reg[45][12]  ( .ip(n16119), .ck(clk), .q(\x[45][12] ) );
  dp_1 \x_reg[45][11]  ( .ip(n16118), .ck(clk), .q(\x[45][11] ) );
  dp_1 \x_reg[45][10]  ( .ip(n16117), .ck(clk), .q(\x[45][10] ) );
  dp_1 \x_reg[45][9]  ( .ip(n16116), .ck(clk), .q(\x[45][9] ) );
  dp_1 \x_reg[45][8]  ( .ip(n16115), .ck(clk), .q(\x[45][8] ) );
  dp_1 \x_reg[45][7]  ( .ip(n16114), .ck(clk), .q(\x[45][7] ) );
  dp_1 \x_reg[45][6]  ( .ip(n16113), .ck(clk), .q(\x[45][6] ) );
  dp_1 \x_reg[45][5]  ( .ip(n16112), .ck(clk), .q(\x[45][5] ) );
  dp_1 \x_reg[45][4]  ( .ip(n16111), .ck(clk), .q(\x[45][4] ) );
  dp_1 \x_reg[45][3]  ( .ip(n16110), .ck(clk), .q(\x[45][3] ) );
  dp_1 \x_reg[45][2]  ( .ip(n16109), .ck(clk), .q(\x[45][2] ) );
  dp_1 \x_reg[45][1]  ( .ip(n16108), .ck(clk), .q(\x[45][1] ) );
  dp_1 \x_reg[45][0]  ( .ip(n16107), .ck(clk), .q(\x[45][0] ) );
  dp_1 \x_reg[44][15]  ( .ip(n16106), .ck(clk), .q(\x[44][15] ) );
  dp_1 \x_reg[44][14]  ( .ip(n16105), .ck(clk), .q(\x[44][14] ) );
  dp_1 \x_reg[44][13]  ( .ip(n16104), .ck(clk), .q(\x[44][13] ) );
  dp_1 \x_reg[44][12]  ( .ip(n16103), .ck(clk), .q(\x[44][12] ) );
  dp_1 \x_reg[44][11]  ( .ip(n16102), .ck(clk), .q(\x[44][11] ) );
  dp_1 \x_reg[44][10]  ( .ip(n16101), .ck(clk), .q(\x[44][10] ) );
  dp_1 \x_reg[44][9]  ( .ip(n16100), .ck(clk), .q(\x[44][9] ) );
  dp_1 \x_reg[44][8]  ( .ip(n16099), .ck(clk), .q(\x[44][8] ) );
  dp_1 \x_reg[44][7]  ( .ip(n16098), .ck(clk), .q(\x[44][7] ) );
  dp_1 \x_reg[44][6]  ( .ip(n16097), .ck(clk), .q(\x[44][6] ) );
  dp_1 \x_reg[44][5]  ( .ip(n16096), .ck(clk), .q(\x[44][5] ) );
  dp_1 \x_reg[44][4]  ( .ip(n16095), .ck(clk), .q(\x[44][4] ) );
  dp_1 \x_reg[44][3]  ( .ip(n16094), .ck(clk), .q(\x[44][3] ) );
  dp_1 \x_reg[44][2]  ( .ip(n16093), .ck(clk), .q(\x[44][2] ) );
  dp_1 \x_reg[44][1]  ( .ip(n16092), .ck(clk), .q(\x[44][1] ) );
  dp_1 \x_reg[44][0]  ( .ip(n16091), .ck(clk), .q(\x[44][0] ) );
  dp_1 \x_reg[43][15]  ( .ip(n16090), .ck(clk), .q(\x[43][15] ) );
  dp_1 \x_reg[43][14]  ( .ip(n16089), .ck(clk), .q(\x[43][14] ) );
  dp_1 \x_reg[43][13]  ( .ip(n16088), .ck(clk), .q(\x[43][13] ) );
  dp_1 \x_reg[43][12]  ( .ip(n16087), .ck(clk), .q(\x[43][12] ) );
  dp_1 \x_reg[43][11]  ( .ip(n16086), .ck(clk), .q(\x[43][11] ) );
  dp_1 \x_reg[43][10]  ( .ip(n16085), .ck(clk), .q(\x[43][10] ) );
  dp_1 \x_reg[43][9]  ( .ip(n16084), .ck(clk), .q(\x[43][9] ) );
  dp_1 \x_reg[43][8]  ( .ip(n16083), .ck(clk), .q(\x[43][8] ) );
  dp_1 \x_reg[43][7]  ( .ip(n16082), .ck(clk), .q(\x[43][7] ) );
  dp_1 \x_reg[43][6]  ( .ip(n16081), .ck(clk), .q(\x[43][6] ) );
  dp_1 \x_reg[43][5]  ( .ip(n16080), .ck(clk), .q(\x[43][5] ) );
  dp_1 \x_reg[43][4]  ( .ip(n16079), .ck(clk), .q(\x[43][4] ) );
  dp_1 \x_reg[43][3]  ( .ip(n16078), .ck(clk), .q(\x[43][3] ) );
  dp_1 \x_reg[43][2]  ( .ip(n16077), .ck(clk), .q(\x[43][2] ) );
  dp_1 \x_reg[43][1]  ( .ip(n16076), .ck(clk), .q(\x[43][1] ) );
  dp_1 \x_reg[43][0]  ( .ip(n16075), .ck(clk), .q(\x[43][0] ) );
  dp_1 \x_reg[42][15]  ( .ip(n16074), .ck(clk), .q(\x[42][15] ) );
  dp_1 \x_reg[42][14]  ( .ip(n16073), .ck(clk), .q(\x[42][14] ) );
  dp_1 \x_reg[42][13]  ( .ip(n16072), .ck(clk), .q(\x[42][13] ) );
  dp_1 \x_reg[42][12]  ( .ip(n16071), .ck(clk), .q(\x[42][12] ) );
  dp_1 \x_reg[42][11]  ( .ip(n16070), .ck(clk), .q(\x[42][11] ) );
  dp_1 \x_reg[42][10]  ( .ip(n16069), .ck(clk), .q(\x[42][10] ) );
  dp_1 \x_reg[42][9]  ( .ip(n16068), .ck(clk), .q(\x[42][9] ) );
  dp_1 \x_reg[42][8]  ( .ip(n16067), .ck(clk), .q(\x[42][8] ) );
  dp_1 \x_reg[42][7]  ( .ip(n16066), .ck(clk), .q(\x[42][7] ) );
  dp_1 \x_reg[42][6]  ( .ip(n16065), .ck(clk), .q(\x[42][6] ) );
  dp_1 \x_reg[42][5]  ( .ip(n16064), .ck(clk), .q(\x[42][5] ) );
  dp_1 \x_reg[42][4]  ( .ip(n16063), .ck(clk), .q(\x[42][4] ) );
  dp_1 \x_reg[42][3]  ( .ip(n16062), .ck(clk), .q(\x[42][3] ) );
  dp_1 \x_reg[42][2]  ( .ip(n16061), .ck(clk), .q(\x[42][2] ) );
  dp_1 \x_reg[42][1]  ( .ip(n16060), .ck(clk), .q(\x[42][1] ) );
  dp_1 \x_reg[42][0]  ( .ip(n16059), .ck(clk), .q(\x[42][0] ) );
  dp_1 \x_reg[41][15]  ( .ip(n16058), .ck(clk), .q(\x[41][15] ) );
  dp_1 \x_reg[41][14]  ( .ip(n16057), .ck(clk), .q(\x[41][14] ) );
  dp_1 \x_reg[41][13]  ( .ip(n16056), .ck(clk), .q(\x[41][13] ) );
  dp_1 \x_reg[41][12]  ( .ip(n16055), .ck(clk), .q(\x[41][12] ) );
  dp_1 \x_reg[41][11]  ( .ip(n16054), .ck(clk), .q(\x[41][11] ) );
  dp_1 \x_reg[41][10]  ( .ip(n16053), .ck(clk), .q(\x[41][10] ) );
  dp_1 \x_reg[41][9]  ( .ip(n16052), .ck(clk), .q(\x[41][9] ) );
  dp_1 \x_reg[41][8]  ( .ip(n16051), .ck(clk), .q(\x[41][8] ) );
  dp_1 \x_reg[41][7]  ( .ip(n16050), .ck(clk), .q(\x[41][7] ) );
  dp_1 \x_reg[41][6]  ( .ip(n16049), .ck(clk), .q(\x[41][6] ) );
  dp_1 \x_reg[41][5]  ( .ip(n16048), .ck(clk), .q(\x[41][5] ) );
  dp_1 \x_reg[41][4]  ( .ip(n16047), .ck(clk), .q(\x[41][4] ) );
  dp_1 \x_reg[41][3]  ( .ip(n16046), .ck(clk), .q(\x[41][3] ) );
  dp_1 \x_reg[41][2]  ( .ip(n16045), .ck(clk), .q(\x[41][2] ) );
  dp_1 \x_reg[41][1]  ( .ip(n16044), .ck(clk), .q(\x[41][1] ) );
  dp_1 \x_reg[41][0]  ( .ip(n16043), .ck(clk), .q(\x[41][0] ) );
  dp_1 \x_reg[40][15]  ( .ip(n16042), .ck(clk), .q(\x[40][15] ) );
  dp_1 \x_reg[40][14]  ( .ip(n16041), .ck(clk), .q(\x[40][14] ) );
  dp_1 \x_reg[40][13]  ( .ip(n16040), .ck(clk), .q(\x[40][13] ) );
  dp_1 \x_reg[40][12]  ( .ip(n16039), .ck(clk), .q(\x[40][12] ) );
  dp_1 \x_reg[40][11]  ( .ip(n16038), .ck(clk), .q(\x[40][11] ) );
  dp_1 \x_reg[40][10]  ( .ip(n16037), .ck(clk), .q(\x[40][10] ) );
  dp_1 \x_reg[40][9]  ( .ip(n16036), .ck(clk), .q(\x[40][9] ) );
  dp_1 \x_reg[40][8]  ( .ip(n16035), .ck(clk), .q(\x[40][8] ) );
  dp_1 \x_reg[40][7]  ( .ip(n16034), .ck(clk), .q(\x[40][7] ) );
  dp_1 \x_reg[40][6]  ( .ip(n16033), .ck(clk), .q(\x[40][6] ) );
  dp_1 \x_reg[40][5]  ( .ip(n16032), .ck(clk), .q(\x[40][5] ) );
  dp_1 \x_reg[40][4]  ( .ip(n16031), .ck(clk), .q(\x[40][4] ) );
  dp_1 \x_reg[40][3]  ( .ip(n16030), .ck(clk), .q(\x[40][3] ) );
  dp_1 \x_reg[40][2]  ( .ip(n16029), .ck(clk), .q(\x[40][2] ) );
  dp_1 \x_reg[40][1]  ( .ip(n16028), .ck(clk), .q(\x[40][1] ) );
  dp_1 \x_reg[40][0]  ( .ip(n16027), .ck(clk), .q(\x[40][0] ) );
  dp_1 \x_reg[39][15]  ( .ip(n16026), .ck(clk), .q(\x[39][15] ) );
  dp_1 \x_reg[39][14]  ( .ip(n16025), .ck(clk), .q(\x[39][14] ) );
  dp_1 \x_reg[39][13]  ( .ip(n16024), .ck(clk), .q(\x[39][13] ) );
  dp_1 \x_reg[39][12]  ( .ip(n16023), .ck(clk), .q(\x[39][12] ) );
  dp_1 \x_reg[39][11]  ( .ip(n16022), .ck(clk), .q(\x[39][11] ) );
  dp_1 \x_reg[39][10]  ( .ip(n16021), .ck(clk), .q(\x[39][10] ) );
  dp_1 \x_reg[39][9]  ( .ip(n16020), .ck(clk), .q(\x[39][9] ) );
  dp_1 \x_reg[39][8]  ( .ip(n16019), .ck(clk), .q(\x[39][8] ) );
  dp_1 \x_reg[39][7]  ( .ip(n16018), .ck(clk), .q(\x[39][7] ) );
  dp_1 \x_reg[39][6]  ( .ip(n16017), .ck(clk), .q(\x[39][6] ) );
  dp_1 \x_reg[39][5]  ( .ip(n16016), .ck(clk), .q(\x[39][5] ) );
  dp_1 \x_reg[39][4]  ( .ip(n16015), .ck(clk), .q(\x[39][4] ) );
  dp_1 \x_reg[39][3]  ( .ip(n16014), .ck(clk), .q(\x[39][3] ) );
  dp_1 \x_reg[39][2]  ( .ip(n16013), .ck(clk), .q(\x[39][2] ) );
  dp_1 \x_reg[39][1]  ( .ip(n16012), .ck(clk), .q(\x[39][1] ) );
  dp_1 \x_reg[39][0]  ( .ip(n16011), .ck(clk), .q(\x[39][0] ) );
  dp_1 \x_reg[38][15]  ( .ip(n16010), .ck(clk), .q(\x[38][15] ) );
  dp_1 \x_reg[38][14]  ( .ip(n16009), .ck(clk), .q(\x[38][14] ) );
  dp_1 \x_reg[38][13]  ( .ip(n16008), .ck(clk), .q(\x[38][13] ) );
  dp_1 \x_reg[38][12]  ( .ip(n16007), .ck(clk), .q(\x[38][12] ) );
  dp_1 \x_reg[38][11]  ( .ip(n16006), .ck(clk), .q(\x[38][11] ) );
  dp_1 \x_reg[38][10]  ( .ip(n16005), .ck(clk), .q(\x[38][10] ) );
  dp_1 \x_reg[38][9]  ( .ip(n16004), .ck(clk), .q(\x[38][9] ) );
  dp_1 \x_reg[38][8]  ( .ip(n16003), .ck(clk), .q(\x[38][8] ) );
  dp_1 \x_reg[38][7]  ( .ip(n16002), .ck(clk), .q(\x[38][7] ) );
  dp_1 \x_reg[38][6]  ( .ip(n16001), .ck(clk), .q(\x[38][6] ) );
  dp_1 \x_reg[38][5]  ( .ip(n16000), .ck(clk), .q(\x[38][5] ) );
  dp_1 \x_reg[38][4]  ( .ip(n15999), .ck(clk), .q(\x[38][4] ) );
  dp_1 \x_reg[38][3]  ( .ip(n15998), .ck(clk), .q(\x[38][3] ) );
  dp_1 \x_reg[38][2]  ( .ip(n15997), .ck(clk), .q(\x[38][2] ) );
  dp_1 \x_reg[38][1]  ( .ip(n15996), .ck(clk), .q(\x[38][1] ) );
  dp_1 \x_reg[38][0]  ( .ip(n15995), .ck(clk), .q(\x[38][0] ) );
  dp_1 \x_reg[37][15]  ( .ip(n15994), .ck(clk), .q(\x[37][15] ) );
  dp_1 \x_reg[37][14]  ( .ip(n15993), .ck(clk), .q(\x[37][14] ) );
  dp_1 \x_reg[37][13]  ( .ip(n15992), .ck(clk), .q(\x[37][13] ) );
  dp_1 \x_reg[37][12]  ( .ip(n15991), .ck(clk), .q(\x[37][12] ) );
  dp_1 \x_reg[37][11]  ( .ip(n15990), .ck(clk), .q(\x[37][11] ) );
  dp_1 \x_reg[37][10]  ( .ip(n15989), .ck(clk), .q(\x[37][10] ) );
  dp_1 \x_reg[37][9]  ( .ip(n15988), .ck(clk), .q(\x[37][9] ) );
  dp_1 \x_reg[37][8]  ( .ip(n15987), .ck(clk), .q(\x[37][8] ) );
  dp_1 \x_reg[37][7]  ( .ip(n15986), .ck(clk), .q(\x[37][7] ) );
  dp_1 \x_reg[37][6]  ( .ip(n15985), .ck(clk), .q(\x[37][6] ) );
  dp_1 \x_reg[37][5]  ( .ip(n15984), .ck(clk), .q(\x[37][5] ) );
  dp_1 \x_reg[37][4]  ( .ip(n15983), .ck(clk), .q(\x[37][4] ) );
  dp_1 \x_reg[37][3]  ( .ip(n15982), .ck(clk), .q(\x[37][3] ) );
  dp_1 \x_reg[37][2]  ( .ip(n15981), .ck(clk), .q(\x[37][2] ) );
  dp_1 \x_reg[37][1]  ( .ip(n15980), .ck(clk), .q(\x[37][1] ) );
  dp_1 \x_reg[37][0]  ( .ip(n15979), .ck(clk), .q(\x[37][0] ) );
  dp_1 \x_reg[36][15]  ( .ip(n15978), .ck(clk), .q(\x[36][15] ) );
  dp_1 \x_reg[36][14]  ( .ip(n15977), .ck(clk), .q(\x[36][14] ) );
  dp_1 \x_reg[36][13]  ( .ip(n15976), .ck(clk), .q(\x[36][13] ) );
  dp_1 \x_reg[36][12]  ( .ip(n15975), .ck(clk), .q(\x[36][12] ) );
  dp_1 \x_reg[36][11]  ( .ip(n15974), .ck(clk), .q(\x[36][11] ) );
  dp_1 \x_reg[36][10]  ( .ip(n15973), .ck(clk), .q(\x[36][10] ) );
  dp_1 \x_reg[36][9]  ( .ip(n15972), .ck(clk), .q(\x[36][9] ) );
  dp_1 \x_reg[36][8]  ( .ip(n15971), .ck(clk), .q(\x[36][8] ) );
  dp_1 \x_reg[36][7]  ( .ip(n15970), .ck(clk), .q(\x[36][7] ) );
  dp_1 \x_reg[36][6]  ( .ip(n15969), .ck(clk), .q(\x[36][6] ) );
  dp_1 \x_reg[36][5]  ( .ip(n15968), .ck(clk), .q(\x[36][5] ) );
  dp_1 \x_reg[36][4]  ( .ip(n15967), .ck(clk), .q(\x[36][4] ) );
  dp_1 \x_reg[36][3]  ( .ip(n15966), .ck(clk), .q(\x[36][3] ) );
  dp_1 \x_reg[36][2]  ( .ip(n15965), .ck(clk), .q(\x[36][2] ) );
  dp_1 \x_reg[36][1]  ( .ip(n15964), .ck(clk), .q(\x[36][1] ) );
  dp_1 \x_reg[36][0]  ( .ip(n15963), .ck(clk), .q(\x[36][0] ) );
  dp_1 \x_reg[35][15]  ( .ip(n15962), .ck(clk), .q(\x[35][15] ) );
  dp_1 \x_reg[35][14]  ( .ip(n15961), .ck(clk), .q(\x[35][14] ) );
  dp_1 \x_reg[35][13]  ( .ip(n15960), .ck(clk), .q(\x[35][13] ) );
  dp_1 \x_reg[35][12]  ( .ip(n15959), .ck(clk), .q(\x[35][12] ) );
  dp_1 \x_reg[35][11]  ( .ip(n15958), .ck(clk), .q(\x[35][11] ) );
  dp_1 \x_reg[35][10]  ( .ip(n15957), .ck(clk), .q(\x[35][10] ) );
  dp_1 \x_reg[35][9]  ( .ip(n15956), .ck(clk), .q(\x[35][9] ) );
  dp_1 \x_reg[35][8]  ( .ip(n15955), .ck(clk), .q(\x[35][8] ) );
  dp_1 \x_reg[35][7]  ( .ip(n15954), .ck(clk), .q(\x[35][7] ) );
  dp_1 \x_reg[35][6]  ( .ip(n15953), .ck(clk), .q(\x[35][6] ) );
  dp_1 \x_reg[35][5]  ( .ip(n15952), .ck(clk), .q(\x[35][5] ) );
  dp_1 \x_reg[35][4]  ( .ip(n15951), .ck(clk), .q(\x[35][4] ) );
  dp_1 \x_reg[35][3]  ( .ip(n15950), .ck(clk), .q(\x[35][3] ) );
  dp_1 \x_reg[35][2]  ( .ip(n15949), .ck(clk), .q(\x[35][2] ) );
  dp_1 \x_reg[35][1]  ( .ip(n15948), .ck(clk), .q(\x[35][1] ) );
  dp_1 \x_reg[35][0]  ( .ip(n15947), .ck(clk), .q(\x[35][0] ) );
  dp_1 \x_reg[34][15]  ( .ip(n15946), .ck(clk), .q(\x[34][15] ) );
  dp_1 \x_reg[34][14]  ( .ip(n15945), .ck(clk), .q(\x[34][14] ) );
  dp_1 \x_reg[34][13]  ( .ip(n15944), .ck(clk), .q(\x[34][13] ) );
  dp_1 \x_reg[34][12]  ( .ip(n15943), .ck(clk), .q(\x[34][12] ) );
  dp_1 \x_reg[34][11]  ( .ip(n15942), .ck(clk), .q(\x[34][11] ) );
  dp_1 \x_reg[34][10]  ( .ip(n15941), .ck(clk), .q(\x[34][10] ) );
  dp_1 \x_reg[34][9]  ( .ip(n15940), .ck(clk), .q(\x[34][9] ) );
  dp_1 \x_reg[34][8]  ( .ip(n15939), .ck(clk), .q(\x[34][8] ) );
  dp_1 \x_reg[34][7]  ( .ip(n15938), .ck(clk), .q(\x[34][7] ) );
  dp_1 \x_reg[34][6]  ( .ip(n15937), .ck(clk), .q(\x[34][6] ) );
  dp_1 \x_reg[34][5]  ( .ip(n15936), .ck(clk), .q(\x[34][5] ) );
  dp_1 \x_reg[34][4]  ( .ip(n15935), .ck(clk), .q(\x[34][4] ) );
  dp_1 \x_reg[34][3]  ( .ip(n15934), .ck(clk), .q(\x[34][3] ) );
  dp_1 \x_reg[34][2]  ( .ip(n15933), .ck(clk), .q(\x[34][2] ) );
  dp_1 \x_reg[34][1]  ( .ip(n15932), .ck(clk), .q(\x[34][1] ) );
  dp_1 \x_reg[34][0]  ( .ip(n15931), .ck(clk), .q(\x[34][0] ) );
  dp_1 \x_reg[33][15]  ( .ip(n15930), .ck(clk), .q(\x[33][15] ) );
  dp_1 \x_reg[33][14]  ( .ip(n15929), .ck(clk), .q(\x[33][14] ) );
  dp_1 \x_reg[33][13]  ( .ip(n15928), .ck(clk), .q(\x[33][13] ) );
  dp_1 \x_reg[33][12]  ( .ip(n15927), .ck(clk), .q(\x[33][12] ) );
  dp_1 \x_reg[33][11]  ( .ip(n15926), .ck(clk), .q(\x[33][11] ) );
  dp_1 \x_reg[33][10]  ( .ip(n15925), .ck(clk), .q(\x[33][10] ) );
  dp_1 \x_reg[33][9]  ( .ip(n15924), .ck(clk), .q(\x[33][9] ) );
  dp_1 \x_reg[33][8]  ( .ip(n15923), .ck(clk), .q(\x[33][8] ) );
  dp_1 \x_reg[33][7]  ( .ip(n15922), .ck(clk), .q(\x[33][7] ) );
  dp_1 \x_reg[33][6]  ( .ip(n15921), .ck(clk), .q(\x[33][6] ) );
  dp_1 \x_reg[33][5]  ( .ip(n15920), .ck(clk), .q(\x[33][5] ) );
  dp_1 \x_reg[33][4]  ( .ip(n15919), .ck(clk), .q(\x[33][4] ) );
  dp_1 \x_reg[33][3]  ( .ip(n15918), .ck(clk), .q(\x[33][3] ) );
  dp_1 \x_reg[33][2]  ( .ip(n15917), .ck(clk), .q(\x[33][2] ) );
  dp_1 \x_reg[33][1]  ( .ip(n15916), .ck(clk), .q(\x[33][1] ) );
  dp_1 \x_reg[33][0]  ( .ip(n15915), .ck(clk), .q(\x[33][0] ) );
  dp_1 \x_reg[32][15]  ( .ip(n15914), .ck(clk), .q(\x[32][15] ) );
  dp_1 \x_reg[32][14]  ( .ip(n15913), .ck(clk), .q(\x[32][14] ) );
  dp_1 \x_reg[32][13]  ( .ip(n15912), .ck(clk), .q(\x[32][13] ) );
  dp_1 \x_reg[32][12]  ( .ip(n15911), .ck(clk), .q(\x[32][12] ) );
  dp_1 \x_reg[32][11]  ( .ip(n15910), .ck(clk), .q(\x[32][11] ) );
  dp_1 \x_reg[32][10]  ( .ip(n15909), .ck(clk), .q(\x[32][10] ) );
  dp_1 \x_reg[32][9]  ( .ip(n15908), .ck(clk), .q(\x[32][9] ) );
  dp_1 \x_reg[32][8]  ( .ip(n15907), .ck(clk), .q(\x[32][8] ) );
  dp_1 \x_reg[32][7]  ( .ip(n15906), .ck(clk), .q(\x[32][7] ) );
  dp_1 \x_reg[32][6]  ( .ip(n15905), .ck(clk), .q(\x[32][6] ) );
  dp_1 \x_reg[32][5]  ( .ip(n15904), .ck(clk), .q(\x[32][5] ) );
  dp_1 \x_reg[32][4]  ( .ip(n15903), .ck(clk), .q(\x[32][4] ) );
  dp_1 \x_reg[32][3]  ( .ip(n15902), .ck(clk), .q(\x[32][3] ) );
  dp_1 \x_reg[32][2]  ( .ip(n15901), .ck(clk), .q(\x[32][2] ) );
  dp_1 \x_reg[32][1]  ( .ip(n15900), .ck(clk), .q(\x[32][1] ) );
  dp_1 \x_reg[32][0]  ( .ip(n15899), .ck(clk), .q(\x[32][0] ) );
  dp_1 \x_reg[31][15]  ( .ip(n15898), .ck(clk), .q(\x[31][15] ) );
  dp_1 \x_reg[31][14]  ( .ip(n15897), .ck(clk), .q(\x[31][14] ) );
  dp_1 \x_reg[31][13]  ( .ip(n15896), .ck(clk), .q(\x[31][13] ) );
  dp_1 \x_reg[31][12]  ( .ip(n15895), .ck(clk), .q(\x[31][12] ) );
  dp_1 \x_reg[31][11]  ( .ip(n15894), .ck(clk), .q(\x[31][11] ) );
  dp_1 \x_reg[31][10]  ( .ip(n15893), .ck(clk), .q(\x[31][10] ) );
  dp_1 \x_reg[31][9]  ( .ip(n15892), .ck(clk), .q(\x[31][9] ) );
  dp_1 \x_reg[31][8]  ( .ip(n15891), .ck(clk), .q(\x[31][8] ) );
  dp_1 \x_reg[31][7]  ( .ip(n15890), .ck(clk), .q(\x[31][7] ) );
  dp_1 \x_reg[31][6]  ( .ip(n15889), .ck(clk), .q(\x[31][6] ) );
  dp_1 \x_reg[31][5]  ( .ip(n15888), .ck(clk), .q(\x[31][5] ) );
  dp_1 \x_reg[31][4]  ( .ip(n15887), .ck(clk), .q(\x[31][4] ) );
  dp_1 \x_reg[31][3]  ( .ip(n15886), .ck(clk), .q(\x[31][3] ) );
  dp_1 \x_reg[31][2]  ( .ip(n15885), .ck(clk), .q(\x[31][2] ) );
  dp_1 \x_reg[31][1]  ( .ip(n15884), .ck(clk), .q(\x[31][1] ) );
  dp_1 \x_reg[31][0]  ( .ip(n15883), .ck(clk), .q(\x[31][0] ) );
  dp_1 \x_reg[30][15]  ( .ip(n15882), .ck(clk), .q(\x[30][15] ) );
  dp_1 \x_reg[30][14]  ( .ip(n15881), .ck(clk), .q(\x[30][14] ) );
  dp_1 \x_reg[30][13]  ( .ip(n15880), .ck(clk), .q(\x[30][13] ) );
  dp_1 \x_reg[30][12]  ( .ip(n15879), .ck(clk), .q(\x[30][12] ) );
  dp_1 \x_reg[30][11]  ( .ip(n15878), .ck(clk), .q(\x[30][11] ) );
  dp_1 \x_reg[30][10]  ( .ip(n15877), .ck(clk), .q(\x[30][10] ) );
  dp_1 \x_reg[30][9]  ( .ip(n15876), .ck(clk), .q(\x[30][9] ) );
  dp_1 \x_reg[30][8]  ( .ip(n15875), .ck(clk), .q(\x[30][8] ) );
  dp_1 \x_reg[30][7]  ( .ip(n15874), .ck(clk), .q(\x[30][7] ) );
  dp_1 \x_reg[30][6]  ( .ip(n15873), .ck(clk), .q(\x[30][6] ) );
  dp_1 \x_reg[30][5]  ( .ip(n15872), .ck(clk), .q(\x[30][5] ) );
  dp_1 \x_reg[30][4]  ( .ip(n15871), .ck(clk), .q(\x[30][4] ) );
  dp_1 \x_reg[30][3]  ( .ip(n15870), .ck(clk), .q(\x[30][3] ) );
  dp_1 \x_reg[30][2]  ( .ip(n15869), .ck(clk), .q(\x[30][2] ) );
  dp_1 \x_reg[30][1]  ( .ip(n15868), .ck(clk), .q(\x[30][1] ) );
  dp_1 \x_reg[30][0]  ( .ip(n15867), .ck(clk), .q(\x[30][0] ) );
  dp_1 \x_reg[29][15]  ( .ip(n15866), .ck(clk), .q(\x[29][15] ) );
  dp_1 \x_reg[29][14]  ( .ip(n15865), .ck(clk), .q(\x[29][14] ) );
  dp_1 \x_reg[29][13]  ( .ip(n15864), .ck(clk), .q(\x[29][13] ) );
  dp_1 \x_reg[29][12]  ( .ip(n15863), .ck(clk), .q(\x[29][12] ) );
  dp_1 \x_reg[29][11]  ( .ip(n15862), .ck(clk), .q(\x[29][11] ) );
  dp_1 \x_reg[29][10]  ( .ip(n15861), .ck(clk), .q(\x[29][10] ) );
  dp_1 \x_reg[29][9]  ( .ip(n15860), .ck(clk), .q(\x[29][9] ) );
  dp_1 \x_reg[29][8]  ( .ip(n15859), .ck(clk), .q(\x[29][8] ) );
  dp_1 \x_reg[29][7]  ( .ip(n15858), .ck(clk), .q(\x[29][7] ) );
  dp_1 \x_reg[29][6]  ( .ip(n15857), .ck(clk), .q(\x[29][6] ) );
  dp_1 \x_reg[29][5]  ( .ip(n15856), .ck(clk), .q(\x[29][5] ) );
  dp_1 \x_reg[29][4]  ( .ip(n15855), .ck(clk), .q(\x[29][4] ) );
  dp_1 \x_reg[29][3]  ( .ip(n15854), .ck(clk), .q(\x[29][3] ) );
  dp_1 \x_reg[29][2]  ( .ip(n15853), .ck(clk), .q(\x[29][2] ) );
  dp_1 \x_reg[29][1]  ( .ip(n15852), .ck(clk), .q(\x[29][1] ) );
  dp_1 \x_reg[29][0]  ( .ip(n15851), .ck(clk), .q(\x[29][0] ) );
  dp_1 \x_reg[28][15]  ( .ip(n15850), .ck(clk), .q(\x[28][15] ) );
  dp_1 \x_reg[28][14]  ( .ip(n15849), .ck(clk), .q(\x[28][14] ) );
  dp_1 \x_reg[28][13]  ( .ip(n15848), .ck(clk), .q(\x[28][13] ) );
  dp_1 \x_reg[28][12]  ( .ip(n15847), .ck(clk), .q(\x[28][12] ) );
  dp_1 \x_reg[28][11]  ( .ip(n15846), .ck(clk), .q(\x[28][11] ) );
  dp_1 \x_reg[28][10]  ( .ip(n15845), .ck(clk), .q(\x[28][10] ) );
  dp_1 \x_reg[28][9]  ( .ip(n15844), .ck(clk), .q(\x[28][9] ) );
  dp_1 \x_reg[28][8]  ( .ip(n15843), .ck(clk), .q(\x[28][8] ) );
  dp_1 \x_reg[28][7]  ( .ip(n15842), .ck(clk), .q(\x[28][7] ) );
  dp_1 \x_reg[28][6]  ( .ip(n15841), .ck(clk), .q(\x[28][6] ) );
  dp_1 \x_reg[28][5]  ( .ip(n15840), .ck(clk), .q(\x[28][5] ) );
  dp_1 \x_reg[28][4]  ( .ip(n15839), .ck(clk), .q(\x[28][4] ) );
  dp_1 \x_reg[28][3]  ( .ip(n15838), .ck(clk), .q(\x[28][3] ) );
  dp_1 \x_reg[28][2]  ( .ip(n15837), .ck(clk), .q(\x[28][2] ) );
  dp_1 \x_reg[28][1]  ( .ip(n15836), .ck(clk), .q(\x[28][1] ) );
  dp_1 \x_reg[28][0]  ( .ip(n15835), .ck(clk), .q(\x[28][0] ) );
  dp_1 \x_reg[27][15]  ( .ip(n15834), .ck(clk), .q(\x[27][15] ) );
  dp_1 \x_reg[27][14]  ( .ip(n15833), .ck(clk), .q(\x[27][14] ) );
  dp_1 \x_reg[27][13]  ( .ip(n15832), .ck(clk), .q(\x[27][13] ) );
  dp_1 \x_reg[27][12]  ( .ip(n15831), .ck(clk), .q(\x[27][12] ) );
  dp_1 \x_reg[27][11]  ( .ip(n15830), .ck(clk), .q(\x[27][11] ) );
  dp_1 \x_reg[27][10]  ( .ip(n15829), .ck(clk), .q(\x[27][10] ) );
  dp_1 \x_reg[27][9]  ( .ip(n15828), .ck(clk), .q(\x[27][9] ) );
  dp_1 \x_reg[27][8]  ( .ip(n15827), .ck(clk), .q(\x[27][8] ) );
  dp_1 \x_reg[27][7]  ( .ip(n15826), .ck(clk), .q(\x[27][7] ) );
  dp_1 \x_reg[27][6]  ( .ip(n15825), .ck(clk), .q(\x[27][6] ) );
  dp_1 \x_reg[27][5]  ( .ip(n15824), .ck(clk), .q(\x[27][5] ) );
  dp_1 \x_reg[27][4]  ( .ip(n15823), .ck(clk), .q(\x[27][4] ) );
  dp_1 \x_reg[27][3]  ( .ip(n15822), .ck(clk), .q(\x[27][3] ) );
  dp_1 \x_reg[27][2]  ( .ip(n15821), .ck(clk), .q(\x[27][2] ) );
  dp_1 \x_reg[27][1]  ( .ip(n15820), .ck(clk), .q(\x[27][1] ) );
  dp_1 \x_reg[27][0]  ( .ip(n15819), .ck(clk), .q(\x[27][0] ) );
  dp_1 \x_reg[26][15]  ( .ip(n15818), .ck(clk), .q(\x[26][15] ) );
  dp_1 \x_reg[26][14]  ( .ip(n15817), .ck(clk), .q(\x[26][14] ) );
  dp_1 \x_reg[26][13]  ( .ip(n15816), .ck(clk), .q(\x[26][13] ) );
  dp_1 \x_reg[26][12]  ( .ip(n15815), .ck(clk), .q(\x[26][12] ) );
  dp_1 \x_reg[26][11]  ( .ip(n15814), .ck(clk), .q(\x[26][11] ) );
  dp_1 \x_reg[26][10]  ( .ip(n15813), .ck(clk), .q(\x[26][10] ) );
  dp_1 \x_reg[26][9]  ( .ip(n15812), .ck(clk), .q(\x[26][9] ) );
  dp_1 \x_reg[26][8]  ( .ip(n15811), .ck(clk), .q(\x[26][8] ) );
  dp_1 \x_reg[26][7]  ( .ip(n15810), .ck(clk), .q(\x[26][7] ) );
  dp_1 \x_reg[26][6]  ( .ip(n15809), .ck(clk), .q(\x[26][6] ) );
  dp_1 \x_reg[26][5]  ( .ip(n15808), .ck(clk), .q(\x[26][5] ) );
  dp_1 \x_reg[26][4]  ( .ip(n15807), .ck(clk), .q(\x[26][4] ) );
  dp_1 \x_reg[26][3]  ( .ip(n15806), .ck(clk), .q(\x[26][3] ) );
  dp_1 \x_reg[26][2]  ( .ip(n15805), .ck(clk), .q(\x[26][2] ) );
  dp_1 \x_reg[26][1]  ( .ip(n15804), .ck(clk), .q(\x[26][1] ) );
  dp_1 \x_reg[26][0]  ( .ip(n15803), .ck(clk), .q(\x[26][0] ) );
  dp_1 \x_reg[25][15]  ( .ip(n15802), .ck(clk), .q(\x[25][15] ) );
  dp_1 \x_reg[25][14]  ( .ip(n15801), .ck(clk), .q(\x[25][14] ) );
  dp_1 \x_reg[25][13]  ( .ip(n15800), .ck(clk), .q(\x[25][13] ) );
  dp_1 \x_reg[25][12]  ( .ip(n15799), .ck(clk), .q(\x[25][12] ) );
  dp_1 \x_reg[25][11]  ( .ip(n15798), .ck(clk), .q(\x[25][11] ) );
  dp_1 \x_reg[25][10]  ( .ip(n15797), .ck(clk), .q(\x[25][10] ) );
  dp_1 \x_reg[25][9]  ( .ip(n15796), .ck(clk), .q(\x[25][9] ) );
  dp_1 \x_reg[25][8]  ( .ip(n15795), .ck(clk), .q(\x[25][8] ) );
  dp_1 \x_reg[25][7]  ( .ip(n15794), .ck(clk), .q(\x[25][7] ) );
  dp_1 \x_reg[25][6]  ( .ip(n15793), .ck(clk), .q(\x[25][6] ) );
  dp_1 \x_reg[25][5]  ( .ip(n15792), .ck(clk), .q(\x[25][5] ) );
  dp_1 \x_reg[25][4]  ( .ip(n15791), .ck(clk), .q(\x[25][4] ) );
  dp_1 \x_reg[25][3]  ( .ip(n15790), .ck(clk), .q(\x[25][3] ) );
  dp_1 \x_reg[25][2]  ( .ip(n15789), .ck(clk), .q(\x[25][2] ) );
  dp_1 \x_reg[25][1]  ( .ip(n15788), .ck(clk), .q(\x[25][1] ) );
  dp_1 \x_reg[25][0]  ( .ip(n15787), .ck(clk), .q(\x[25][0] ) );
  dp_1 \x_reg[24][15]  ( .ip(n15786), .ck(clk), .q(\x[24][15] ) );
  dp_1 \x_reg[24][14]  ( .ip(n15785), .ck(clk), .q(\x[24][14] ) );
  dp_1 \x_reg[24][13]  ( .ip(n15784), .ck(clk), .q(\x[24][13] ) );
  dp_1 \x_reg[24][12]  ( .ip(n15783), .ck(clk), .q(\x[24][12] ) );
  dp_1 \x_reg[24][11]  ( .ip(n15782), .ck(clk), .q(\x[24][11] ) );
  dp_1 \x_reg[24][10]  ( .ip(n15781), .ck(clk), .q(\x[24][10] ) );
  dp_1 \x_reg[24][9]  ( .ip(n15780), .ck(clk), .q(\x[24][9] ) );
  dp_1 \x_reg[24][8]  ( .ip(n15779), .ck(clk), .q(\x[24][8] ) );
  dp_1 \x_reg[24][7]  ( .ip(n15778), .ck(clk), .q(\x[24][7] ) );
  dp_1 \x_reg[24][6]  ( .ip(n15777), .ck(clk), .q(\x[24][6] ) );
  dp_1 \x_reg[24][5]  ( .ip(n15776), .ck(clk), .q(\x[24][5] ) );
  dp_1 \x_reg[24][4]  ( .ip(n15775), .ck(clk), .q(\x[24][4] ) );
  dp_1 \x_reg[24][3]  ( .ip(n15774), .ck(clk), .q(\x[24][3] ) );
  dp_1 \x_reg[24][2]  ( .ip(n15773), .ck(clk), .q(\x[24][2] ) );
  dp_1 \x_reg[24][1]  ( .ip(n15772), .ck(clk), .q(\x[24][1] ) );
  dp_1 \x_reg[24][0]  ( .ip(n15771), .ck(clk), .q(\x[24][0] ) );
  dp_1 \x_reg[23][15]  ( .ip(n15770), .ck(clk), .q(\x[23][15] ) );
  dp_1 \x_reg[23][14]  ( .ip(n15769), .ck(clk), .q(\x[23][14] ) );
  dp_1 \x_reg[23][13]  ( .ip(n15768), .ck(clk), .q(\x[23][13] ) );
  dp_1 \x_reg[23][12]  ( .ip(n15767), .ck(clk), .q(\x[23][12] ) );
  dp_1 \x_reg[23][11]  ( .ip(n15766), .ck(clk), .q(\x[23][11] ) );
  dp_1 \x_reg[23][10]  ( .ip(n15765), .ck(clk), .q(\x[23][10] ) );
  dp_1 \x_reg[23][9]  ( .ip(n15764), .ck(clk), .q(\x[23][9] ) );
  dp_1 \x_reg[23][8]  ( .ip(n15763), .ck(clk), .q(\x[23][8] ) );
  dp_1 \x_reg[23][7]  ( .ip(n15762), .ck(clk), .q(\x[23][7] ) );
  dp_1 \x_reg[23][6]  ( .ip(n15761), .ck(clk), .q(\x[23][6] ) );
  dp_1 \x_reg[23][5]  ( .ip(n15760), .ck(clk), .q(\x[23][5] ) );
  dp_1 \x_reg[23][4]  ( .ip(n15759), .ck(clk), .q(\x[23][4] ) );
  dp_1 \x_reg[23][3]  ( .ip(n15758), .ck(clk), .q(\x[23][3] ) );
  dp_1 \x_reg[23][2]  ( .ip(n15757), .ck(clk), .q(\x[23][2] ) );
  dp_1 \x_reg[23][1]  ( .ip(n15756), .ck(clk), .q(\x[23][1] ) );
  dp_1 \x_reg[23][0]  ( .ip(n15755), .ck(clk), .q(\x[23][0] ) );
  dp_1 \x_reg[22][15]  ( .ip(n15754), .ck(clk), .q(\x[22][15] ) );
  dp_1 \x_reg[22][14]  ( .ip(n15753), .ck(clk), .q(\x[22][14] ) );
  dp_1 \x_reg[22][13]  ( .ip(n15752), .ck(clk), .q(\x[22][13] ) );
  dp_1 \x_reg[22][12]  ( .ip(n15751), .ck(clk), .q(\x[22][12] ) );
  dp_1 \x_reg[22][11]  ( .ip(n15750), .ck(clk), .q(\x[22][11] ) );
  dp_1 \x_reg[22][10]  ( .ip(n15749), .ck(clk), .q(\x[22][10] ) );
  dp_1 \x_reg[22][9]  ( .ip(n15748), .ck(clk), .q(\x[22][9] ) );
  dp_1 \x_reg[22][8]  ( .ip(n15747), .ck(clk), .q(\x[22][8] ) );
  dp_1 \x_reg[22][7]  ( .ip(n15746), .ck(clk), .q(\x[22][7] ) );
  dp_1 \x_reg[22][6]  ( .ip(n15745), .ck(clk), .q(\x[22][6] ) );
  dp_1 \x_reg[22][5]  ( .ip(n15744), .ck(clk), .q(\x[22][5] ) );
  dp_1 \x_reg[22][4]  ( .ip(n15743), .ck(clk), .q(\x[22][4] ) );
  dp_1 \x_reg[22][3]  ( .ip(n15742), .ck(clk), .q(\x[22][3] ) );
  dp_1 \x_reg[22][2]  ( .ip(n15741), .ck(clk), .q(\x[22][2] ) );
  dp_1 \x_reg[22][1]  ( .ip(n15740), .ck(clk), .q(\x[22][1] ) );
  dp_1 \x_reg[22][0]  ( .ip(n15739), .ck(clk), .q(\x[22][0] ) );
  dp_1 \x_reg[21][15]  ( .ip(n15738), .ck(clk), .q(\x[21][15] ) );
  dp_1 \x_reg[21][14]  ( .ip(n15737), .ck(clk), .q(\x[21][14] ) );
  dp_1 \x_reg[21][13]  ( .ip(n15736), .ck(clk), .q(\x[21][13] ) );
  dp_1 \x_reg[21][12]  ( .ip(n15735), .ck(clk), .q(\x[21][12] ) );
  dp_1 \x_reg[21][11]  ( .ip(n15734), .ck(clk), .q(\x[21][11] ) );
  dp_1 \x_reg[21][10]  ( .ip(n15733), .ck(clk), .q(\x[21][10] ) );
  dp_1 \x_reg[21][9]  ( .ip(n15732), .ck(clk), .q(\x[21][9] ) );
  dp_1 \x_reg[21][8]  ( .ip(n15731), .ck(clk), .q(\x[21][8] ) );
  dp_1 \x_reg[21][7]  ( .ip(n15730), .ck(clk), .q(\x[21][7] ) );
  dp_1 \x_reg[21][6]  ( .ip(n15729), .ck(clk), .q(\x[21][6] ) );
  dp_1 \x_reg[21][5]  ( .ip(n15728), .ck(clk), .q(\x[21][5] ) );
  dp_1 \x_reg[21][4]  ( .ip(n15727), .ck(clk), .q(\x[21][4] ) );
  dp_1 \x_reg[21][3]  ( .ip(n15726), .ck(clk), .q(\x[21][3] ) );
  dp_1 \x_reg[21][2]  ( .ip(n15725), .ck(clk), .q(\x[21][2] ) );
  dp_1 \x_reg[21][1]  ( .ip(n15724), .ck(clk), .q(\x[21][1] ) );
  dp_1 \x_reg[21][0]  ( .ip(n15723), .ck(clk), .q(\x[21][0] ) );
  dp_1 \x_reg[20][15]  ( .ip(n15722), .ck(clk), .q(\x[20][15] ) );
  dp_1 \x_reg[20][14]  ( .ip(n15721), .ck(clk), .q(\x[20][14] ) );
  dp_1 \x_reg[20][13]  ( .ip(n15720), .ck(clk), .q(\x[20][13] ) );
  dp_1 \x_reg[20][12]  ( .ip(n15719), .ck(clk), .q(\x[20][12] ) );
  dp_1 \x_reg[20][11]  ( .ip(n15718), .ck(clk), .q(\x[20][11] ) );
  dp_1 \x_reg[20][10]  ( .ip(n15717), .ck(clk), .q(\x[20][10] ) );
  dp_1 \x_reg[20][9]  ( .ip(n15716), .ck(clk), .q(\x[20][9] ) );
  dp_1 \x_reg[20][8]  ( .ip(n15715), .ck(clk), .q(\x[20][8] ) );
  dp_1 \x_reg[20][7]  ( .ip(n15714), .ck(clk), .q(\x[20][7] ) );
  dp_1 \x_reg[20][6]  ( .ip(n15713), .ck(clk), .q(\x[20][6] ) );
  dp_1 \x_reg[20][5]  ( .ip(n15712), .ck(clk), .q(\x[20][5] ) );
  dp_1 \x_reg[20][4]  ( .ip(n15711), .ck(clk), .q(\x[20][4] ) );
  dp_1 \x_reg[20][3]  ( .ip(n15710), .ck(clk), .q(\x[20][3] ) );
  dp_1 \x_reg[20][2]  ( .ip(n15709), .ck(clk), .q(\x[20][2] ) );
  dp_1 \x_reg[20][1]  ( .ip(n15708), .ck(clk), .q(\x[20][1] ) );
  dp_1 \x_reg[20][0]  ( .ip(n15707), .ck(clk), .q(\x[20][0] ) );
  dp_1 \x_reg[19][15]  ( .ip(n15706), .ck(clk), .q(\x[19][15] ) );
  dp_1 \x_reg[19][14]  ( .ip(n15705), .ck(clk), .q(\x[19][14] ) );
  dp_1 \x_reg[19][13]  ( .ip(n15704), .ck(clk), .q(\x[19][13] ) );
  dp_1 \x_reg[19][12]  ( .ip(n15703), .ck(clk), .q(\x[19][12] ) );
  dp_1 \x_reg[19][11]  ( .ip(n15702), .ck(clk), .q(\x[19][11] ) );
  dp_1 \x_reg[19][10]  ( .ip(n15701), .ck(clk), .q(\x[19][10] ) );
  dp_1 \x_reg[19][9]  ( .ip(n15700), .ck(clk), .q(\x[19][9] ) );
  dp_1 \x_reg[19][8]  ( .ip(n15699), .ck(clk), .q(\x[19][8] ) );
  dp_1 \x_reg[19][7]  ( .ip(n15698), .ck(clk), .q(\x[19][7] ) );
  dp_1 \x_reg[19][6]  ( .ip(n15697), .ck(clk), .q(\x[19][6] ) );
  dp_1 \x_reg[19][5]  ( .ip(n15696), .ck(clk), .q(\x[19][5] ) );
  dp_1 \x_reg[19][4]  ( .ip(n15695), .ck(clk), .q(\x[19][4] ) );
  dp_1 \x_reg[19][3]  ( .ip(n15694), .ck(clk), .q(\x[19][3] ) );
  dp_1 \x_reg[19][2]  ( .ip(n15693), .ck(clk), .q(\x[19][2] ) );
  dp_1 \x_reg[19][1]  ( .ip(n15692), .ck(clk), .q(\x[19][1] ) );
  dp_1 \x_reg[19][0]  ( .ip(n15691), .ck(clk), .q(\x[19][0] ) );
  dp_1 \x_reg[18][15]  ( .ip(n15690), .ck(clk), .q(\x[18][15] ) );
  dp_1 \x_reg[18][14]  ( .ip(n15689), .ck(clk), .q(\x[18][14] ) );
  dp_1 \x_reg[18][13]  ( .ip(n15688), .ck(clk), .q(\x[18][13] ) );
  dp_1 \x_reg[18][12]  ( .ip(n15687), .ck(clk), .q(\x[18][12] ) );
  dp_1 \x_reg[18][11]  ( .ip(n15686), .ck(clk), .q(\x[18][11] ) );
  dp_1 \x_reg[18][10]  ( .ip(n15685), .ck(clk), .q(\x[18][10] ) );
  dp_1 \x_reg[18][9]  ( .ip(n15684), .ck(clk), .q(\x[18][9] ) );
  dp_1 \x_reg[18][8]  ( .ip(n15683), .ck(clk), .q(\x[18][8] ) );
  dp_1 \x_reg[18][7]  ( .ip(n15682), .ck(clk), .q(\x[18][7] ) );
  dp_1 \x_reg[18][6]  ( .ip(n15681), .ck(clk), .q(\x[18][6] ) );
  dp_1 \x_reg[18][5]  ( .ip(n15680), .ck(clk), .q(\x[18][5] ) );
  dp_1 \x_reg[18][4]  ( .ip(n15679), .ck(clk), .q(\x[18][4] ) );
  dp_1 \x_reg[18][3]  ( .ip(n15678), .ck(clk), .q(\x[18][3] ) );
  dp_1 \x_reg[18][2]  ( .ip(n15677), .ck(clk), .q(\x[18][2] ) );
  dp_1 \x_reg[18][1]  ( .ip(n15676), .ck(clk), .q(\x[18][1] ) );
  dp_1 \x_reg[18][0]  ( .ip(n15675), .ck(clk), .q(\x[18][0] ) );
  dp_1 \x_reg[17][15]  ( .ip(n15674), .ck(clk), .q(\x[17][15] ) );
  dp_1 \x_reg[17][14]  ( .ip(n15673), .ck(clk), .q(\x[17][14] ) );
  dp_1 \x_reg[17][13]  ( .ip(n15672), .ck(clk), .q(\x[17][13] ) );
  dp_1 \x_reg[17][12]  ( .ip(n15671), .ck(clk), .q(\x[17][12] ) );
  dp_1 \x_reg[17][11]  ( .ip(n15670), .ck(clk), .q(\x[17][11] ) );
  dp_1 \x_reg[17][10]  ( .ip(n15669), .ck(clk), .q(\x[17][10] ) );
  dp_1 \x_reg[17][9]  ( .ip(n15668), .ck(clk), .q(\x[17][9] ) );
  dp_1 \x_reg[17][8]  ( .ip(n15667), .ck(clk), .q(\x[17][8] ) );
  dp_1 \x_reg[17][7]  ( .ip(n15666), .ck(clk), .q(\x[17][7] ) );
  dp_1 \x_reg[17][6]  ( .ip(n15665), .ck(clk), .q(\x[17][6] ) );
  dp_1 \x_reg[17][5]  ( .ip(n15664), .ck(clk), .q(\x[17][5] ) );
  dp_1 \x_reg[17][4]  ( .ip(n15663), .ck(clk), .q(\x[17][4] ) );
  dp_1 \x_reg[17][3]  ( .ip(n15662), .ck(clk), .q(\x[17][3] ) );
  dp_1 \x_reg[17][2]  ( .ip(n15661), .ck(clk), .q(\x[17][2] ) );
  dp_1 \x_reg[17][1]  ( .ip(n15660), .ck(clk), .q(\x[17][1] ) );
  dp_1 \x_reg[17][0]  ( .ip(n15659), .ck(clk), .q(\x[17][0] ) );
  dp_1 \x_reg[16][15]  ( .ip(n15658), .ck(clk), .q(\x[16][15] ) );
  dp_1 \x_reg[16][14]  ( .ip(n15657), .ck(clk), .q(\x[16][14] ) );
  dp_1 \x_reg[16][13]  ( .ip(n15656), .ck(clk), .q(\x[16][13] ) );
  dp_1 \x_reg[16][12]  ( .ip(n15655), .ck(clk), .q(\x[16][12] ) );
  dp_1 \x_reg[16][11]  ( .ip(n15654), .ck(clk), .q(\x[16][11] ) );
  dp_1 \x_reg[16][10]  ( .ip(n15653), .ck(clk), .q(\x[16][10] ) );
  dp_1 \x_reg[16][9]  ( .ip(n15652), .ck(clk), .q(\x[16][9] ) );
  dp_1 \x_reg[16][8]  ( .ip(n15651), .ck(clk), .q(\x[16][8] ) );
  dp_1 \x_reg[16][7]  ( .ip(n15650), .ck(clk), .q(\x[16][7] ) );
  dp_1 \x_reg[16][6]  ( .ip(n15649), .ck(clk), .q(\x[16][6] ) );
  dp_1 \x_reg[16][5]  ( .ip(n15648), .ck(clk), .q(\x[16][5] ) );
  dp_1 \x_reg[16][4]  ( .ip(n15647), .ck(clk), .q(\x[16][4] ) );
  dp_1 \x_reg[16][3]  ( .ip(n15646), .ck(clk), .q(\x[16][3] ) );
  dp_1 \x_reg[16][2]  ( .ip(n15645), .ck(clk), .q(\x[16][2] ) );
  dp_1 \x_reg[16][1]  ( .ip(n15644), .ck(clk), .q(\x[16][1] ) );
  dp_1 \x_reg[16][0]  ( .ip(n15643), .ck(clk), .q(\x[16][0] ) );
  dp_1 \x_reg[15][15]  ( .ip(n15642), .ck(clk), .q(\x[15][15] ) );
  dp_1 \x_reg[15][14]  ( .ip(n15641), .ck(clk), .q(\x[15][14] ) );
  dp_1 \x_reg[15][13]  ( .ip(n15640), .ck(clk), .q(\x[15][13] ) );
  dp_1 \x_reg[15][12]  ( .ip(n15639), .ck(clk), .q(\x[15][12] ) );
  dp_1 \x_reg[15][11]  ( .ip(n15638), .ck(clk), .q(\x[15][11] ) );
  dp_1 \x_reg[15][10]  ( .ip(n15637), .ck(clk), .q(\x[15][10] ) );
  dp_1 \x_reg[15][9]  ( .ip(n15636), .ck(clk), .q(\x[15][9] ) );
  dp_1 \x_reg[15][8]  ( .ip(n15635), .ck(clk), .q(\x[15][8] ) );
  dp_1 \x_reg[15][7]  ( .ip(n15634), .ck(clk), .q(\x[15][7] ) );
  dp_1 \x_reg[15][6]  ( .ip(n15633), .ck(clk), .q(\x[15][6] ) );
  dp_1 \x_reg[15][5]  ( .ip(n15632), .ck(clk), .q(\x[15][5] ) );
  dp_1 \x_reg[15][4]  ( .ip(n15631), .ck(clk), .q(\x[15][4] ) );
  dp_1 \x_reg[15][3]  ( .ip(n15630), .ck(clk), .q(\x[15][3] ) );
  dp_1 \x_reg[15][2]  ( .ip(n15629), .ck(clk), .q(\x[15][2] ) );
  dp_1 \x_reg[15][1]  ( .ip(n15628), .ck(clk), .q(\x[15][1] ) );
  dp_1 \x_reg[15][0]  ( .ip(n15627), .ck(clk), .q(\x[15][0] ) );
  dp_1 \x_reg[14][15]  ( .ip(n15626), .ck(clk), .q(\x[14][15] ) );
  dp_1 \x_reg[14][14]  ( .ip(n15625), .ck(clk), .q(\x[14][14] ) );
  dp_1 \x_reg[14][13]  ( .ip(n15624), .ck(clk), .q(\x[14][13] ) );
  dp_1 \x_reg[14][12]  ( .ip(n15623), .ck(clk), .q(\x[14][12] ) );
  dp_1 \x_reg[14][11]  ( .ip(n15622), .ck(clk), .q(\x[14][11] ) );
  dp_1 \x_reg[14][10]  ( .ip(n15621), .ck(clk), .q(\x[14][10] ) );
  dp_1 \x_reg[14][9]  ( .ip(n15620), .ck(clk), .q(\x[14][9] ) );
  dp_1 \x_reg[14][8]  ( .ip(n15619), .ck(clk), .q(\x[14][8] ) );
  dp_1 \x_reg[14][7]  ( .ip(n15618), .ck(clk), .q(\x[14][7] ) );
  dp_1 \x_reg[14][6]  ( .ip(n15617), .ck(clk), .q(\x[14][6] ) );
  dp_1 \x_reg[14][5]  ( .ip(n15616), .ck(clk), .q(\x[14][5] ) );
  dp_1 \x_reg[14][4]  ( .ip(n15615), .ck(clk), .q(\x[14][4] ) );
  dp_1 \x_reg[14][3]  ( .ip(n15614), .ck(clk), .q(\x[14][3] ) );
  dp_1 \x_reg[14][2]  ( .ip(n15613), .ck(clk), .q(\x[14][2] ) );
  dp_1 \x_reg[14][1]  ( .ip(n15612), .ck(clk), .q(\x[14][1] ) );
  dp_1 \x_reg[14][0]  ( .ip(n15611), .ck(clk), .q(\x[14][0] ) );
  dp_1 \x_reg[13][15]  ( .ip(n15610), .ck(clk), .q(\x[13][15] ) );
  dp_1 \x_reg[13][14]  ( .ip(n15609), .ck(clk), .q(\x[13][14] ) );
  dp_1 \x_reg[13][13]  ( .ip(n15608), .ck(clk), .q(\x[13][13] ) );
  dp_1 \x_reg[13][12]  ( .ip(n15607), .ck(clk), .q(\x[13][12] ) );
  dp_1 \x_reg[13][11]  ( .ip(n15606), .ck(clk), .q(\x[13][11] ) );
  dp_1 \x_reg[13][10]  ( .ip(n15605), .ck(clk), .q(\x[13][10] ) );
  dp_1 \x_reg[13][9]  ( .ip(n15604), .ck(clk), .q(\x[13][9] ) );
  dp_1 \x_reg[13][8]  ( .ip(n15603), .ck(clk), .q(\x[13][8] ) );
  dp_1 \x_reg[13][7]  ( .ip(n15602), .ck(clk), .q(\x[13][7] ) );
  dp_1 \x_reg[13][6]  ( .ip(n15601), .ck(clk), .q(\x[13][6] ) );
  dp_1 \x_reg[13][5]  ( .ip(n15600), .ck(clk), .q(\x[13][5] ) );
  dp_1 \x_reg[13][4]  ( .ip(n15599), .ck(clk), .q(\x[13][4] ) );
  dp_1 \x_reg[13][3]  ( .ip(n15598), .ck(clk), .q(\x[13][3] ) );
  dp_1 \x_reg[13][2]  ( .ip(n15597), .ck(clk), .q(\x[13][2] ) );
  dp_1 \x_reg[13][1]  ( .ip(n15596), .ck(clk), .q(\x[13][1] ) );
  dp_1 \x_reg[13][0]  ( .ip(n15595), .ck(clk), .q(\x[13][0] ) );
  dp_1 \x_reg[12][15]  ( .ip(n15594), .ck(clk), .q(\x[12][15] ) );
  dp_1 \x_reg[12][14]  ( .ip(n15593), .ck(clk), .q(\x[12][14] ) );
  dp_1 \x_reg[12][13]  ( .ip(n15592), .ck(clk), .q(\x[12][13] ) );
  dp_1 \x_reg[12][12]  ( .ip(n15591), .ck(clk), .q(\x[12][12] ) );
  dp_1 \x_reg[12][11]  ( .ip(n15590), .ck(clk), .q(\x[12][11] ) );
  dp_1 \x_reg[12][10]  ( .ip(n15589), .ck(clk), .q(\x[12][10] ) );
  dp_1 \x_reg[12][9]  ( .ip(n15588), .ck(clk), .q(\x[12][9] ) );
  dp_1 \x_reg[12][8]  ( .ip(n15587), .ck(clk), .q(\x[12][8] ) );
  dp_1 \x_reg[12][7]  ( .ip(n15586), .ck(clk), .q(\x[12][7] ) );
  dp_1 \x_reg[12][6]  ( .ip(n15585), .ck(clk), .q(\x[12][6] ) );
  dp_1 \x_reg[12][5]  ( .ip(n15584), .ck(clk), .q(\x[12][5] ) );
  dp_1 \x_reg[12][4]  ( .ip(n15583), .ck(clk), .q(\x[12][4] ) );
  dp_1 \x_reg[12][3]  ( .ip(n15582), .ck(clk), .q(\x[12][3] ) );
  dp_1 \x_reg[12][2]  ( .ip(n15581), .ck(clk), .q(\x[12][2] ) );
  dp_1 \x_reg[12][1]  ( .ip(n15580), .ck(clk), .q(\x[12][1] ) );
  dp_1 \x_reg[12][0]  ( .ip(n15579), .ck(clk), .q(\x[12][0] ) );
  dp_1 \x_reg[11][15]  ( .ip(n15578), .ck(clk), .q(\x[11][15] ) );
  dp_1 \x_reg[11][14]  ( .ip(n15577), .ck(clk), .q(\x[11][14] ) );
  dp_1 \x_reg[11][13]  ( .ip(n15576), .ck(clk), .q(\x[11][13] ) );
  dp_1 \x_reg[11][12]  ( .ip(n15575), .ck(clk), .q(\x[11][12] ) );
  dp_1 \x_reg[11][11]  ( .ip(n15574), .ck(clk), .q(\x[11][11] ) );
  dp_1 \x_reg[11][10]  ( .ip(n15573), .ck(clk), .q(\x[11][10] ) );
  dp_1 \x_reg[11][9]  ( .ip(n15572), .ck(clk), .q(\x[11][9] ) );
  dp_1 \x_reg[11][8]  ( .ip(n15571), .ck(clk), .q(\x[11][8] ) );
  dp_1 \x_reg[11][7]  ( .ip(n15570), .ck(clk), .q(\x[11][7] ) );
  dp_1 \x_reg[11][6]  ( .ip(n15569), .ck(clk), .q(\x[11][6] ) );
  dp_1 \x_reg[11][5]  ( .ip(n15568), .ck(clk), .q(\x[11][5] ) );
  dp_1 \x_reg[11][4]  ( .ip(n15567), .ck(clk), .q(\x[11][4] ) );
  dp_1 \x_reg[11][3]  ( .ip(n15566), .ck(clk), .q(\x[11][3] ) );
  dp_1 \x_reg[11][2]  ( .ip(n15565), .ck(clk), .q(\x[11][2] ) );
  dp_1 \x_reg[11][1]  ( .ip(n15564), .ck(clk), .q(\x[11][1] ) );
  dp_1 \x_reg[11][0]  ( .ip(n15563), .ck(clk), .q(\x[11][0] ) );
  dp_1 \x_reg[10][15]  ( .ip(n15562), .ck(clk), .q(\x[10][15] ) );
  dp_1 \x_reg[10][14]  ( .ip(n15561), .ck(clk), .q(\x[10][14] ) );
  dp_1 \x_reg[10][13]  ( .ip(n15560), .ck(clk), .q(\x[10][13] ) );
  dp_1 \x_reg[10][12]  ( .ip(n15559), .ck(clk), .q(\x[10][12] ) );
  dp_1 \x_reg[10][11]  ( .ip(n15558), .ck(clk), .q(\x[10][11] ) );
  dp_1 \x_reg[10][10]  ( .ip(n15557), .ck(clk), .q(\x[10][10] ) );
  dp_1 \x_reg[10][9]  ( .ip(n15556), .ck(clk), .q(\x[10][9] ) );
  dp_1 \x_reg[10][8]  ( .ip(n15555), .ck(clk), .q(\x[10][8] ) );
  dp_1 \x_reg[10][7]  ( .ip(n15554), .ck(clk), .q(\x[10][7] ) );
  dp_1 \x_reg[10][6]  ( .ip(n15553), .ck(clk), .q(\x[10][6] ) );
  dp_1 \x_reg[10][5]  ( .ip(n15552), .ck(clk), .q(\x[10][5] ) );
  dp_1 \x_reg[10][4]  ( .ip(n15551), .ck(clk), .q(\x[10][4] ) );
  dp_1 \x_reg[10][3]  ( .ip(n15550), .ck(clk), .q(\x[10][3] ) );
  dp_1 \x_reg[10][2]  ( .ip(n15549), .ck(clk), .q(\x[10][2] ) );
  dp_1 \x_reg[10][1]  ( .ip(n15548), .ck(clk), .q(\x[10][1] ) );
  dp_1 \x_reg[10][0]  ( .ip(n15547), .ck(clk), .q(\x[10][0] ) );
  dp_1 \x_reg[9][15]  ( .ip(n15546), .ck(clk), .q(\x[9][15] ) );
  dp_1 \x_reg[9][14]  ( .ip(n15545), .ck(clk), .q(\x[9][14] ) );
  dp_1 \x_reg[9][13]  ( .ip(n15544), .ck(clk), .q(\x[9][13] ) );
  dp_1 \x_reg[9][12]  ( .ip(n15543), .ck(clk), .q(\x[9][12] ) );
  dp_1 \x_reg[9][11]  ( .ip(n15542), .ck(clk), .q(\x[9][11] ) );
  dp_1 \x_reg[9][10]  ( .ip(n15541), .ck(clk), .q(\x[9][10] ) );
  dp_1 \x_reg[9][9]  ( .ip(n15540), .ck(clk), .q(\x[9][9] ) );
  dp_1 \x_reg[9][8]  ( .ip(n15539), .ck(clk), .q(\x[9][8] ) );
  dp_1 \x_reg[9][7]  ( .ip(n15538), .ck(clk), .q(\x[9][7] ) );
  dp_1 \x_reg[9][6]  ( .ip(n15537), .ck(clk), .q(\x[9][6] ) );
  dp_1 \x_reg[9][5]  ( .ip(n15536), .ck(clk), .q(\x[9][5] ) );
  dp_1 \x_reg[9][4]  ( .ip(n15535), .ck(clk), .q(\x[9][4] ) );
  dp_1 \x_reg[9][3]  ( .ip(n15534), .ck(clk), .q(\x[9][3] ) );
  dp_1 \x_reg[9][2]  ( .ip(n15533), .ck(clk), .q(\x[9][2] ) );
  dp_1 \x_reg[9][1]  ( .ip(n15532), .ck(clk), .q(\x[9][1] ) );
  dp_1 \x_reg[9][0]  ( .ip(n15531), .ck(clk), .q(\x[9][0] ) );
  dp_1 \x_reg[8][15]  ( .ip(n15530), .ck(clk), .q(\x[8][15] ) );
  dp_1 \x_reg[8][14]  ( .ip(n15529), .ck(clk), .q(\x[8][14] ) );
  dp_1 \x_reg[8][13]  ( .ip(n15528), .ck(clk), .q(\x[8][13] ) );
  dp_1 \x_reg[8][12]  ( .ip(n15527), .ck(clk), .q(\x[8][12] ) );
  dp_1 \x_reg[8][11]  ( .ip(n15526), .ck(clk), .q(\x[8][11] ) );
  dp_1 \x_reg[8][10]  ( .ip(n15525), .ck(clk), .q(\x[8][10] ) );
  dp_1 \x_reg[8][9]  ( .ip(n15524), .ck(clk), .q(\x[8][9] ) );
  dp_1 \x_reg[8][8]  ( .ip(n15523), .ck(clk), .q(\x[8][8] ) );
  dp_1 \x_reg[8][7]  ( .ip(n15522), .ck(clk), .q(\x[8][7] ) );
  dp_1 \x_reg[8][6]  ( .ip(n15521), .ck(clk), .q(\x[8][6] ) );
  dp_1 \x_reg[8][5]  ( .ip(n15520), .ck(clk), .q(\x[8][5] ) );
  dp_1 \x_reg[8][4]  ( .ip(n15519), .ck(clk), .q(\x[8][4] ) );
  dp_1 \x_reg[8][3]  ( .ip(n15518), .ck(clk), .q(\x[8][3] ) );
  dp_1 \x_reg[8][2]  ( .ip(n15517), .ck(clk), .q(\x[8][2] ) );
  dp_1 \x_reg[8][1]  ( .ip(n15516), .ck(clk), .q(\x[8][1] ) );
  dp_1 \x_reg[8][0]  ( .ip(n15515), .ck(clk), .q(\x[8][0] ) );
  dp_1 \x_reg[7][15]  ( .ip(n15514), .ck(clk), .q(\x[7][15] ) );
  dp_1 \x_reg[7][14]  ( .ip(n15513), .ck(clk), .q(\x[7][14] ) );
  dp_1 \x_reg[7][13]  ( .ip(n15512), .ck(clk), .q(\x[7][13] ) );
  dp_1 \x_reg[7][12]  ( .ip(n15511), .ck(clk), .q(\x[7][12] ) );
  dp_1 \x_reg[7][11]  ( .ip(n15510), .ck(clk), .q(\x[7][11] ) );
  dp_1 \x_reg[7][10]  ( .ip(n15509), .ck(clk), .q(\x[7][10] ) );
  dp_1 \x_reg[7][9]  ( .ip(n15508), .ck(clk), .q(\x[7][9] ) );
  dp_1 \x_reg[7][8]  ( .ip(n15507), .ck(clk), .q(\x[7][8] ) );
  dp_1 \x_reg[7][7]  ( .ip(n15506), .ck(clk), .q(\x[7][7] ) );
  dp_1 \x_reg[7][6]  ( .ip(n15505), .ck(clk), .q(\x[7][6] ) );
  dp_1 \x_reg[7][5]  ( .ip(n15504), .ck(clk), .q(\x[7][5] ) );
  dp_1 \x_reg[7][4]  ( .ip(n15503), .ck(clk), .q(\x[7][4] ) );
  dp_1 \x_reg[7][3]  ( .ip(n15502), .ck(clk), .q(\x[7][3] ) );
  dp_1 \x_reg[7][2]  ( .ip(n15501), .ck(clk), .q(\x[7][2] ) );
  dp_1 \x_reg[7][1]  ( .ip(n15500), .ck(clk), .q(\x[7][1] ) );
  dp_1 \x_reg[7][0]  ( .ip(n15499), .ck(clk), .q(\x[7][0] ) );
  dp_1 \x_reg[6][15]  ( .ip(n15498), .ck(clk), .q(\x[6][15] ) );
  dp_1 \x_reg[6][14]  ( .ip(n15497), .ck(clk), .q(\x[6][14] ) );
  dp_1 \x_reg[6][13]  ( .ip(n15496), .ck(clk), .q(\x[6][13] ) );
  dp_1 \x_reg[6][12]  ( .ip(n15495), .ck(clk), .q(\x[6][12] ) );
  dp_1 \x_reg[6][11]  ( .ip(n15494), .ck(clk), .q(\x[6][11] ) );
  dp_1 \x_reg[6][10]  ( .ip(n15493), .ck(clk), .q(\x[6][10] ) );
  dp_1 \x_reg[6][9]  ( .ip(n15492), .ck(clk), .q(\x[6][9] ) );
  dp_1 \x_reg[6][8]  ( .ip(n15491), .ck(clk), .q(\x[6][8] ) );
  dp_1 \x_reg[6][7]  ( .ip(n15490), .ck(clk), .q(\x[6][7] ) );
  dp_1 \x_reg[6][6]  ( .ip(n15489), .ck(clk), .q(\x[6][6] ) );
  dp_1 \x_reg[6][5]  ( .ip(n15488), .ck(clk), .q(\x[6][5] ) );
  dp_1 \x_reg[6][4]  ( .ip(n15487), .ck(clk), .q(\x[6][4] ) );
  dp_1 \x_reg[6][3]  ( .ip(n15486), .ck(clk), .q(\x[6][3] ) );
  dp_1 \x_reg[6][2]  ( .ip(n15485), .ck(clk), .q(\x[6][2] ) );
  dp_1 \x_reg[6][1]  ( .ip(n15484), .ck(clk), .q(\x[6][1] ) );
  dp_1 \x_reg[6][0]  ( .ip(n15483), .ck(clk), .q(\x[6][0] ) );
  dp_1 \x_reg[5][15]  ( .ip(n15482), .ck(clk), .q(\x[5][15] ) );
  dp_1 \x_reg[5][14]  ( .ip(n15481), .ck(clk), .q(\x[5][14] ) );
  dp_1 \x_reg[5][13]  ( .ip(n15480), .ck(clk), .q(\x[5][13] ) );
  dp_1 \x_reg[5][12]  ( .ip(n15479), .ck(clk), .q(\x[5][12] ) );
  dp_1 \x_reg[5][11]  ( .ip(n15478), .ck(clk), .q(\x[5][11] ) );
  dp_1 \x_reg[5][10]  ( .ip(n15477), .ck(clk), .q(\x[5][10] ) );
  dp_1 \x_reg[5][9]  ( .ip(n15476), .ck(clk), .q(\x[5][9] ) );
  dp_1 \x_reg[5][8]  ( .ip(n15475), .ck(clk), .q(\x[5][8] ) );
  dp_1 \x_reg[5][7]  ( .ip(n15474), .ck(clk), .q(\x[5][7] ) );
  dp_1 \x_reg[5][6]  ( .ip(n15473), .ck(clk), .q(\x[5][6] ) );
  dp_1 \x_reg[5][5]  ( .ip(n15472), .ck(clk), .q(\x[5][5] ) );
  dp_1 \x_reg[5][4]  ( .ip(n15471), .ck(clk), .q(\x[5][4] ) );
  dp_1 \x_reg[5][3]  ( .ip(n15470), .ck(clk), .q(\x[5][3] ) );
  dp_1 \x_reg[5][2]  ( .ip(n15469), .ck(clk), .q(\x[5][2] ) );
  dp_1 \x_reg[5][1]  ( .ip(n15468), .ck(clk), .q(\x[5][1] ) );
  dp_1 \x_reg[5][0]  ( .ip(n15467), .ck(clk), .q(\x[5][0] ) );
  dp_1 \x_reg[4][15]  ( .ip(n15466), .ck(clk), .q(\x[4][15] ) );
  dp_1 \x_reg[4][14]  ( .ip(n15465), .ck(clk), .q(\x[4][14] ) );
  dp_1 \x_reg[4][13]  ( .ip(n15464), .ck(clk), .q(\x[4][13] ) );
  dp_1 \x_reg[4][12]  ( .ip(n15463), .ck(clk), .q(\x[4][12] ) );
  dp_1 \x_reg[4][11]  ( .ip(n15462), .ck(clk), .q(\x[4][11] ) );
  dp_1 \x_reg[4][10]  ( .ip(n15461), .ck(clk), .q(\x[4][10] ) );
  dp_1 \x_reg[4][9]  ( .ip(n15460), .ck(clk), .q(\x[4][9] ) );
  dp_1 \x_reg[4][8]  ( .ip(n15459), .ck(clk), .q(\x[4][8] ) );
  dp_1 \x_reg[4][7]  ( .ip(n15458), .ck(clk), .q(\x[4][7] ) );
  dp_1 \x_reg[4][6]  ( .ip(n15457), .ck(clk), .q(\x[4][6] ) );
  dp_1 \x_reg[4][5]  ( .ip(n15456), .ck(clk), .q(\x[4][5] ) );
  dp_1 \x_reg[4][4]  ( .ip(n15455), .ck(clk), .q(\x[4][4] ) );
  dp_1 \x_reg[4][3]  ( .ip(n15454), .ck(clk), .q(\x[4][3] ) );
  dp_1 \x_reg[4][2]  ( .ip(n15453), .ck(clk), .q(\x[4][2] ) );
  dp_1 \x_reg[4][1]  ( .ip(n15452), .ck(clk), .q(\x[4][1] ) );
  dp_1 \x_reg[4][0]  ( .ip(n15451), .ck(clk), .q(\x[4][0] ) );
  dp_1 \x_reg[3][15]  ( .ip(n15450), .ck(clk), .q(\x[3][15] ) );
  dp_1 \x_reg[3][14]  ( .ip(n15449), .ck(clk), .q(\x[3][14] ) );
  dp_1 \x_reg[3][13]  ( .ip(n15448), .ck(clk), .q(\x[3][13] ) );
  dp_1 \x_reg[3][12]  ( .ip(n15447), .ck(clk), .q(\x[3][12] ) );
  dp_1 \x_reg[3][11]  ( .ip(n15446), .ck(clk), .q(\x[3][11] ) );
  dp_1 \x_reg[3][10]  ( .ip(n15445), .ck(clk), .q(\x[3][10] ) );
  dp_1 \x_reg[3][9]  ( .ip(n15444), .ck(clk), .q(\x[3][9] ) );
  dp_1 \x_reg[3][8]  ( .ip(n15443), .ck(clk), .q(\x[3][8] ) );
  dp_1 \x_reg[3][7]  ( .ip(n15442), .ck(clk), .q(\x[3][7] ) );
  dp_1 \x_reg[3][6]  ( .ip(n15441), .ck(clk), .q(\x[3][6] ) );
  dp_1 \x_reg[3][5]  ( .ip(n15440), .ck(clk), .q(\x[3][5] ) );
  dp_1 \x_reg[3][4]  ( .ip(n15439), .ck(clk), .q(\x[3][4] ) );
  dp_1 \x_reg[3][3]  ( .ip(n15438), .ck(clk), .q(\x[3][3] ) );
  dp_1 \x_reg[3][2]  ( .ip(n15437), .ck(clk), .q(\x[3][2] ) );
  dp_1 \x_reg[3][1]  ( .ip(n15436), .ck(clk), .q(\x[3][1] ) );
  dp_1 \x_reg[3][0]  ( .ip(n15435), .ck(clk), .q(\x[3][0] ) );
  dp_1 \x_reg[2][15]  ( .ip(n15434), .ck(clk), .q(\x[2][15] ) );
  dp_1 \x_reg[2][14]  ( .ip(n15433), .ck(clk), .q(\x[2][14] ) );
  dp_1 \x_reg[2][13]  ( .ip(n15432), .ck(clk), .q(\x[2][13] ) );
  dp_1 \x_reg[2][12]  ( .ip(n15431), .ck(clk), .q(\x[2][12] ) );
  dp_1 \x_reg[2][11]  ( .ip(n15430), .ck(clk), .q(\x[2][11] ) );
  dp_1 \x_reg[2][10]  ( .ip(n15429), .ck(clk), .q(\x[2][10] ) );
  dp_1 \x_reg[2][9]  ( .ip(n15428), .ck(clk), .q(\x[2][9] ) );
  dp_1 \x_reg[2][8]  ( .ip(n15427), .ck(clk), .q(\x[2][8] ) );
  dp_1 \x_reg[2][7]  ( .ip(n15426), .ck(clk), .q(\x[2][7] ) );
  dp_1 \x_reg[2][6]  ( .ip(n15425), .ck(clk), .q(\x[2][6] ) );
  dp_1 \x_reg[2][5]  ( .ip(n15424), .ck(clk), .q(\x[2][5] ) );
  dp_1 \x_reg[2][4]  ( .ip(n15423), .ck(clk), .q(\x[2][4] ) );
  dp_1 \x_reg[2][3]  ( .ip(n15422), .ck(clk), .q(\x[2][3] ) );
  dp_1 \x_reg[2][2]  ( .ip(n15421), .ck(clk), .q(\x[2][2] ) );
  dp_1 \x_reg[2][1]  ( .ip(n15420), .ck(clk), .q(\x[2][1] ) );
  dp_1 \x_reg[2][0]  ( .ip(n15419), .ck(clk), .q(\x[2][0] ) );
  dp_1 \x_reg[1][15]  ( .ip(n15418), .ck(clk), .q(\x[1][15] ) );
  dp_1 \x_reg[1][14]  ( .ip(n15417), .ck(clk), .q(\x[1][14] ) );
  dp_1 \x_reg[1][13]  ( .ip(n15416), .ck(clk), .q(\x[1][13] ) );
  dp_1 \x_reg[1][12]  ( .ip(n15415), .ck(clk), .q(\x[1][12] ) );
  dp_1 \x_reg[1][11]  ( .ip(n15414), .ck(clk), .q(\x[1][11] ) );
  dp_1 \x_reg[1][10]  ( .ip(n15413), .ck(clk), .q(\x[1][10] ) );
  dp_1 \x_reg[1][9]  ( .ip(n15412), .ck(clk), .q(\x[1][9] ) );
  dp_1 \x_reg[1][8]  ( .ip(n15411), .ck(clk), .q(\x[1][8] ) );
  dp_1 \x_reg[1][7]  ( .ip(n15410), .ck(clk), .q(\x[1][7] ) );
  dp_1 \x_reg[1][6]  ( .ip(n15409), .ck(clk), .q(\x[1][6] ) );
  dp_1 \x_reg[1][5]  ( .ip(n15408), .ck(clk), .q(\x[1][5] ) );
  dp_1 \x_reg[1][4]  ( .ip(n15407), .ck(clk), .q(\x[1][4] ) );
  dp_1 \x_reg[1][3]  ( .ip(n15406), .ck(clk), .q(\x[1][3] ) );
  dp_1 \x_reg[1][2]  ( .ip(n15405), .ck(clk), .q(\x[1][2] ) );
  dp_1 \x_reg[1][1]  ( .ip(n15404), .ck(clk), .q(\x[1][1] ) );
  dp_1 \x_reg[1][0]  ( .ip(n15403), .ck(clk), .q(\x[1][0] ) );
  dp_1 \x_reg[0][15]  ( .ip(n15402), .ck(clk), .q(\x[0][15] ) );
  dp_1 \x_reg[0][14]  ( .ip(n15401), .ck(clk), .q(\x[0][14] ) );
  dp_1 \x_reg[0][13]  ( .ip(n15400), .ck(clk), .q(\x[0][13] ) );
  dp_1 \x_reg[0][12]  ( .ip(n15399), .ck(clk), .q(\x[0][12] ) );
  dp_1 \x_reg[0][11]  ( .ip(n15398), .ck(clk), .q(\x[0][11] ) );
  dp_1 \x_reg[0][10]  ( .ip(n15397), .ck(clk), .q(\x[0][10] ) );
  dp_1 \x_reg[0][9]  ( .ip(n15396), .ck(clk), .q(\x[0][9] ) );
  dp_1 \x_reg[0][8]  ( .ip(n15395), .ck(clk), .q(\x[0][8] ) );
  dp_1 \x_reg[0][7]  ( .ip(n15394), .ck(clk), .q(\x[0][7] ) );
  dp_1 \x_reg[0][6]  ( .ip(n15393), .ck(clk), .q(\x[0][6] ) );
  dp_1 \x_reg[0][5]  ( .ip(n15392), .ck(clk), .q(\x[0][5] ) );
  dp_1 \x_reg[0][4]  ( .ip(n15391), .ck(clk), .q(\x[0][4] ) );
  dp_1 \x_reg[0][3]  ( .ip(n15390), .ck(clk), .q(\x[0][3] ) );
  dp_1 \x_reg[0][2]  ( .ip(n15389), .ck(clk), .q(\x[0][2] ) );
  dp_1 \x_reg[0][1]  ( .ip(n15388), .ck(clk), .q(\x[0][1] ) );
  dp_1 \x_reg[0][0]  ( .ip(n15387), .ck(clk), .q(\x[0][0] ) );
  dp_1 sig_rdy_reg ( .ip(n15386), .ck(clk), .q(sig_ready) );
  dp_1 \LUT_reg[119][15]  ( .ip(n15385), .ck(clk), .q(\LUT[119][15] ) );
  dp_1 \LUT_reg[119][14]  ( .ip(n15384), .ck(clk), .q(\LUT[119][14] ) );
  dp_1 \LUT_reg[119][13]  ( .ip(n15383), .ck(clk), .q(\LUT[119][13] ) );
  dp_1 \LUT_reg[119][12]  ( .ip(n15382), .ck(clk), .q(\LUT[119][12] ) );
  dp_1 \LUT_reg[119][11]  ( .ip(n15381), .ck(clk), .q(\LUT[119][11] ) );
  dp_1 \LUT_reg[119][10]  ( .ip(n15380), .ck(clk), .q(\LUT[119][10] ) );
  dp_1 \LUT_reg[119][9]  ( .ip(n15379), .ck(clk), .q(\LUT[119][9] ) );
  dp_1 \LUT_reg[119][8]  ( .ip(n15378), .ck(clk), .q(\LUT[119][8] ) );
  dp_1 \LUT_reg[119][7]  ( .ip(n15377), .ck(clk), .q(\LUT[119][7] ) );
  dp_1 \LUT_reg[119][6]  ( .ip(n15376), .ck(clk), .q(\LUT[119][6] ) );
  dp_1 \LUT_reg[119][5]  ( .ip(n15375), .ck(clk), .q(\LUT[119][5] ) );
  dp_1 \LUT_reg[119][4]  ( .ip(n15374), .ck(clk), .q(\LUT[119][4] ) );
  dp_1 \LUT_reg[119][3]  ( .ip(n15373), .ck(clk), .q(\LUT[119][3] ) );
  dp_1 \LUT_reg[119][2]  ( .ip(n15372), .ck(clk), .q(\LUT[119][2] ) );
  dp_1 \LUT_reg[119][1]  ( .ip(n15371), .ck(clk), .q(\LUT[119][1] ) );
  dp_1 \LUT_reg[119][0]  ( .ip(n15370), .ck(clk), .q(\LUT[119][0] ) );
  dp_1 \LUT_reg[118][15]  ( .ip(n15369), .ck(clk), .q(\LUT[118][15] ) );
  dp_1 \LUT_reg[118][14]  ( .ip(n15368), .ck(clk), .q(\LUT[118][14] ) );
  dp_1 \LUT_reg[118][13]  ( .ip(n15367), .ck(clk), .q(\LUT[118][13] ) );
  dp_1 \LUT_reg[118][12]  ( .ip(n15366), .ck(clk), .q(\LUT[118][12] ) );
  dp_1 \LUT_reg[118][11]  ( .ip(n15365), .ck(clk), .q(\LUT[118][11] ) );
  dp_1 \LUT_reg[118][10]  ( .ip(n15364), .ck(clk), .q(\LUT[118][10] ) );
  dp_1 \LUT_reg[118][9]  ( .ip(n15363), .ck(clk), .q(\LUT[118][9] ) );
  dp_1 \LUT_reg[118][8]  ( .ip(n15362), .ck(clk), .q(\LUT[118][8] ) );
  dp_1 \LUT_reg[118][7]  ( .ip(n15361), .ck(clk), .q(\LUT[118][7] ) );
  dp_1 \LUT_reg[118][6]  ( .ip(n15360), .ck(clk), .q(\LUT[118][6] ) );
  dp_1 \LUT_reg[118][5]  ( .ip(n15359), .ck(clk), .q(\LUT[118][5] ) );
  dp_1 \LUT_reg[118][4]  ( .ip(n15358), .ck(clk), .q(\LUT[118][4] ) );
  dp_1 \LUT_reg[118][3]  ( .ip(n15357), .ck(clk), .q(\LUT[118][3] ) );
  dp_1 \LUT_reg[118][2]  ( .ip(n15356), .ck(clk), .q(\LUT[118][2] ) );
  dp_1 \LUT_reg[118][1]  ( .ip(n15355), .ck(clk), .q(\LUT[118][1] ) );
  dp_1 \LUT_reg[118][0]  ( .ip(n15354), .ck(clk), .q(\LUT[118][0] ) );
  dp_1 \LUT_reg[117][15]  ( .ip(n15353), .ck(clk), .q(\LUT[117][15] ) );
  dp_1 \LUT_reg[117][14]  ( .ip(n15352), .ck(clk), .q(\LUT[117][14] ) );
  dp_1 \LUT_reg[117][13]  ( .ip(n15351), .ck(clk), .q(\LUT[117][13] ) );
  dp_1 \LUT_reg[117][12]  ( .ip(n15350), .ck(clk), .q(\LUT[117][12] ) );
  dp_1 \LUT_reg[117][11]  ( .ip(n15349), .ck(clk), .q(\LUT[117][11] ) );
  dp_1 \LUT_reg[117][10]  ( .ip(n15348), .ck(clk), .q(\LUT[117][10] ) );
  dp_1 \LUT_reg[117][9]  ( .ip(n15347), .ck(clk), .q(\LUT[117][9] ) );
  dp_1 \LUT_reg[117][8]  ( .ip(n15346), .ck(clk), .q(\LUT[117][8] ) );
  dp_1 \LUT_reg[117][7]  ( .ip(n15345), .ck(clk), .q(\LUT[117][7] ) );
  dp_1 \LUT_reg[117][6]  ( .ip(n15344), .ck(clk), .q(\LUT[117][6] ) );
  dp_1 \LUT_reg[117][5]  ( .ip(n15343), .ck(clk), .q(\LUT[117][5] ) );
  dp_1 \LUT_reg[117][4]  ( .ip(n15342), .ck(clk), .q(\LUT[117][4] ) );
  dp_1 \LUT_reg[117][3]  ( .ip(n15341), .ck(clk), .q(\LUT[117][3] ) );
  dp_1 \LUT_reg[117][2]  ( .ip(n15340), .ck(clk), .q(\LUT[117][2] ) );
  dp_1 \LUT_reg[117][1]  ( .ip(n15339), .ck(clk), .q(\LUT[117][1] ) );
  dp_1 \LUT_reg[117][0]  ( .ip(n15338), .ck(clk), .q(\LUT[117][0] ) );
  dp_1 \LUT_reg[116][15]  ( .ip(n15337), .ck(clk), .q(\LUT[116][15] ) );
  dp_1 \LUT_reg[116][14]  ( .ip(n15336), .ck(clk), .q(\LUT[116][14] ) );
  dp_1 \LUT_reg[116][13]  ( .ip(n15335), .ck(clk), .q(\LUT[116][13] ) );
  dp_1 \LUT_reg[116][12]  ( .ip(n15334), .ck(clk), .q(\LUT[116][12] ) );
  dp_1 \LUT_reg[116][11]  ( .ip(n15333), .ck(clk), .q(\LUT[116][11] ) );
  dp_1 \LUT_reg[116][10]  ( .ip(n15332), .ck(clk), .q(\LUT[116][10] ) );
  dp_1 \LUT_reg[116][9]  ( .ip(n15331), .ck(clk), .q(\LUT[116][9] ) );
  dp_1 \LUT_reg[116][8]  ( .ip(n15330), .ck(clk), .q(\LUT[116][8] ) );
  dp_1 \LUT_reg[116][7]  ( .ip(n15329), .ck(clk), .q(\LUT[116][7] ) );
  dp_1 \LUT_reg[116][6]  ( .ip(n15328), .ck(clk), .q(\LUT[116][6] ) );
  dp_1 \LUT_reg[116][5]  ( .ip(n15327), .ck(clk), .q(\LUT[116][5] ) );
  dp_1 \LUT_reg[116][4]  ( .ip(n15326), .ck(clk), .q(\LUT[116][4] ) );
  dp_1 \LUT_reg[116][3]  ( .ip(n15325), .ck(clk), .q(\LUT[116][3] ) );
  dp_1 \LUT_reg[116][2]  ( .ip(n15324), .ck(clk), .q(\LUT[116][2] ) );
  dp_1 \LUT_reg[116][1]  ( .ip(n15323), .ck(clk), .q(\LUT[116][1] ) );
  dp_1 \LUT_reg[116][0]  ( .ip(n15322), .ck(clk), .q(\LUT[116][0] ) );
  dp_1 \LUT_reg[115][15]  ( .ip(n15321), .ck(clk), .q(\LUT[115][15] ) );
  dp_1 \LUT_reg[115][14]  ( .ip(n15320), .ck(clk), .q(\LUT[115][14] ) );
  dp_1 \LUT_reg[115][13]  ( .ip(n15319), .ck(clk), .q(\LUT[115][13] ) );
  dp_1 \LUT_reg[115][12]  ( .ip(n15318), .ck(clk), .q(\LUT[115][12] ) );
  dp_1 \LUT_reg[115][11]  ( .ip(n15317), .ck(clk), .q(\LUT[115][11] ) );
  dp_1 \LUT_reg[115][10]  ( .ip(n15316), .ck(clk), .q(\LUT[115][10] ) );
  dp_1 \LUT_reg[115][9]  ( .ip(n15315), .ck(clk), .q(\LUT[115][9] ) );
  dp_1 \LUT_reg[115][8]  ( .ip(n15314), .ck(clk), .q(\LUT[115][8] ) );
  dp_1 \LUT_reg[115][7]  ( .ip(n15313), .ck(clk), .q(\LUT[115][7] ) );
  dp_1 \LUT_reg[115][6]  ( .ip(n15312), .ck(clk), .q(\LUT[115][6] ) );
  dp_1 \LUT_reg[115][5]  ( .ip(n15311), .ck(clk), .q(\LUT[115][5] ) );
  dp_1 \LUT_reg[115][4]  ( .ip(n15310), .ck(clk), .q(\LUT[115][4] ) );
  dp_1 \LUT_reg[115][3]  ( .ip(n15309), .ck(clk), .q(\LUT[115][3] ) );
  dp_1 \LUT_reg[115][2]  ( .ip(n15308), .ck(clk), .q(\LUT[115][2] ) );
  dp_1 \LUT_reg[115][1]  ( .ip(n15307), .ck(clk), .q(\LUT[115][1] ) );
  dp_1 \LUT_reg[115][0]  ( .ip(n15306), .ck(clk), .q(\LUT[115][0] ) );
  dp_1 \LUT_reg[114][15]  ( .ip(n15305), .ck(clk), .q(\LUT[114][15] ) );
  dp_1 \LUT_reg[114][14]  ( .ip(n15304), .ck(clk), .q(\LUT[114][14] ) );
  dp_1 \LUT_reg[114][13]  ( .ip(n15303), .ck(clk), .q(\LUT[114][13] ) );
  dp_1 \LUT_reg[114][12]  ( .ip(n15302), .ck(clk), .q(\LUT[114][12] ) );
  dp_1 \LUT_reg[114][11]  ( .ip(n15301), .ck(clk), .q(\LUT[114][11] ) );
  dp_1 \LUT_reg[114][10]  ( .ip(n15300), .ck(clk), .q(\LUT[114][10] ) );
  dp_1 \LUT_reg[114][9]  ( .ip(n15299), .ck(clk), .q(\LUT[114][9] ) );
  dp_1 \LUT_reg[114][8]  ( .ip(n15298), .ck(clk), .q(\LUT[114][8] ) );
  dp_1 \LUT_reg[114][7]  ( .ip(n15297), .ck(clk), .q(\LUT[114][7] ) );
  dp_1 \LUT_reg[114][6]  ( .ip(n15296), .ck(clk), .q(\LUT[114][6] ) );
  dp_1 \LUT_reg[114][5]  ( .ip(n15295), .ck(clk), .q(\LUT[114][5] ) );
  dp_1 \LUT_reg[114][4]  ( .ip(n15294), .ck(clk), .q(\LUT[114][4] ) );
  dp_1 \LUT_reg[114][3]  ( .ip(n15293), .ck(clk), .q(\LUT[114][3] ) );
  dp_1 \LUT_reg[114][2]  ( .ip(n15292), .ck(clk), .q(\LUT[114][2] ) );
  dp_1 \LUT_reg[114][1]  ( .ip(n15291), .ck(clk), .q(\LUT[114][1] ) );
  dp_1 \LUT_reg[114][0]  ( .ip(n15290), .ck(clk), .q(\LUT[114][0] ) );
  dp_1 \LUT_reg[113][15]  ( .ip(n15289), .ck(clk), .q(\LUT[113][15] ) );
  dp_1 \LUT_reg[113][14]  ( .ip(n15288), .ck(clk), .q(\LUT[113][14] ) );
  dp_1 \LUT_reg[113][13]  ( .ip(n15287), .ck(clk), .q(\LUT[113][13] ) );
  dp_1 \LUT_reg[113][12]  ( .ip(n15286), .ck(clk), .q(\LUT[113][12] ) );
  dp_1 \LUT_reg[113][11]  ( .ip(n15285), .ck(clk), .q(\LUT[113][11] ) );
  dp_1 \LUT_reg[113][10]  ( .ip(n15284), .ck(clk), .q(\LUT[113][10] ) );
  dp_1 \LUT_reg[113][9]  ( .ip(n15283), .ck(clk), .q(\LUT[113][9] ) );
  dp_1 \LUT_reg[113][8]  ( .ip(n15282), .ck(clk), .q(\LUT[113][8] ) );
  dp_1 \LUT_reg[113][7]  ( .ip(n15281), .ck(clk), .q(\LUT[113][7] ) );
  dp_1 \LUT_reg[113][6]  ( .ip(n15280), .ck(clk), .q(\LUT[113][6] ) );
  dp_1 \LUT_reg[113][5]  ( .ip(n15279), .ck(clk), .q(\LUT[113][5] ) );
  dp_1 \LUT_reg[113][4]  ( .ip(n15278), .ck(clk), .q(\LUT[113][4] ) );
  dp_1 \LUT_reg[113][3]  ( .ip(n15277), .ck(clk), .q(\LUT[113][3] ) );
  dp_1 \LUT_reg[113][2]  ( .ip(n15276), .ck(clk), .q(\LUT[113][2] ) );
  dp_1 \LUT_reg[113][1]  ( .ip(n15275), .ck(clk), .q(\LUT[113][1] ) );
  dp_1 \LUT_reg[113][0]  ( .ip(n15274), .ck(clk), .q(\LUT[113][0] ) );
  dp_1 \LUT_reg[112][15]  ( .ip(n15273), .ck(clk), .q(\LUT[112][15] ) );
  dp_1 \LUT_reg[112][14]  ( .ip(n15272), .ck(clk), .q(\LUT[112][14] ) );
  dp_1 \LUT_reg[112][13]  ( .ip(n15271), .ck(clk), .q(\LUT[112][13] ) );
  dp_1 \LUT_reg[112][12]  ( .ip(n15270), .ck(clk), .q(\LUT[112][12] ) );
  dp_1 \LUT_reg[112][11]  ( .ip(n15269), .ck(clk), .q(\LUT[112][11] ) );
  dp_1 \LUT_reg[112][10]  ( .ip(n15268), .ck(clk), .q(\LUT[112][10] ) );
  dp_1 \LUT_reg[112][9]  ( .ip(n15267), .ck(clk), .q(\LUT[112][9] ) );
  dp_1 \LUT_reg[112][8]  ( .ip(n15266), .ck(clk), .q(\LUT[112][8] ) );
  dp_1 \LUT_reg[112][7]  ( .ip(n15265), .ck(clk), .q(\LUT[112][7] ) );
  dp_1 \LUT_reg[112][6]  ( .ip(n15264), .ck(clk), .q(\LUT[112][6] ) );
  dp_1 \LUT_reg[112][5]  ( .ip(n15263), .ck(clk), .q(\LUT[112][5] ) );
  dp_1 \LUT_reg[112][4]  ( .ip(n15262), .ck(clk), .q(\LUT[112][4] ) );
  dp_1 \LUT_reg[112][3]  ( .ip(n15261), .ck(clk), .q(\LUT[112][3] ) );
  dp_1 \LUT_reg[112][2]  ( .ip(n15260), .ck(clk), .q(\LUT[112][2] ) );
  dp_1 \LUT_reg[112][1]  ( .ip(n15259), .ck(clk), .q(\LUT[112][1] ) );
  dp_1 \LUT_reg[112][0]  ( .ip(n15258), .ck(clk), .q(\LUT[112][0] ) );
  dp_1 \LUT_reg[111][15]  ( .ip(n15257), .ck(clk), .q(\LUT[111][15] ) );
  dp_1 \LUT_reg[111][14]  ( .ip(n15256), .ck(clk), .q(\LUT[111][14] ) );
  dp_1 \LUT_reg[111][13]  ( .ip(n15255), .ck(clk), .q(\LUT[111][13] ) );
  dp_1 \LUT_reg[111][12]  ( .ip(n15254), .ck(clk), .q(\LUT[111][12] ) );
  dp_1 \LUT_reg[111][11]  ( .ip(n15253), .ck(clk), .q(\LUT[111][11] ) );
  dp_1 \LUT_reg[111][10]  ( .ip(n15252), .ck(clk), .q(\LUT[111][10] ) );
  dp_1 \LUT_reg[111][9]  ( .ip(n15251), .ck(clk), .q(\LUT[111][9] ) );
  dp_1 \LUT_reg[111][8]  ( .ip(n15250), .ck(clk), .q(\LUT[111][8] ) );
  dp_1 \LUT_reg[111][7]  ( .ip(n15249), .ck(clk), .q(\LUT[111][7] ) );
  dp_1 \LUT_reg[111][6]  ( .ip(n15248), .ck(clk), .q(\LUT[111][6] ) );
  dp_1 \LUT_reg[111][5]  ( .ip(n15247), .ck(clk), .q(\LUT[111][5] ) );
  dp_1 \LUT_reg[111][4]  ( .ip(n15246), .ck(clk), .q(\LUT[111][4] ) );
  dp_1 \LUT_reg[111][3]  ( .ip(n15245), .ck(clk), .q(\LUT[111][3] ) );
  dp_1 \LUT_reg[111][2]  ( .ip(n15244), .ck(clk), .q(\LUT[111][2] ) );
  dp_1 \LUT_reg[111][1]  ( .ip(n15243), .ck(clk), .q(\LUT[111][1] ) );
  dp_1 \LUT_reg[111][0]  ( .ip(n15242), .ck(clk), .q(\LUT[111][0] ) );
  dp_1 \LUT_reg[110][15]  ( .ip(n15241), .ck(clk), .q(\LUT[110][15] ) );
  dp_1 \LUT_reg[110][14]  ( .ip(n15240), .ck(clk), .q(\LUT[110][14] ) );
  dp_1 \LUT_reg[110][13]  ( .ip(n15239), .ck(clk), .q(\LUT[110][13] ) );
  dp_1 \LUT_reg[110][12]  ( .ip(n15238), .ck(clk), .q(\LUT[110][12] ) );
  dp_1 \LUT_reg[110][11]  ( .ip(n15237), .ck(clk), .q(\LUT[110][11] ) );
  dp_1 \LUT_reg[110][10]  ( .ip(n15236), .ck(clk), .q(\LUT[110][10] ) );
  dp_1 \LUT_reg[110][9]  ( .ip(n15235), .ck(clk), .q(\LUT[110][9] ) );
  dp_1 \LUT_reg[110][8]  ( .ip(n15234), .ck(clk), .q(\LUT[110][8] ) );
  dp_1 \LUT_reg[110][7]  ( .ip(n15233), .ck(clk), .q(\LUT[110][7] ) );
  dp_1 \LUT_reg[110][6]  ( .ip(n15232), .ck(clk), .q(\LUT[110][6] ) );
  dp_1 \LUT_reg[110][5]  ( .ip(n15231), .ck(clk), .q(\LUT[110][5] ) );
  dp_1 \LUT_reg[110][4]  ( .ip(n15230), .ck(clk), .q(\LUT[110][4] ) );
  dp_1 \LUT_reg[110][3]  ( .ip(n15229), .ck(clk), .q(\LUT[110][3] ) );
  dp_1 \LUT_reg[110][2]  ( .ip(n15228), .ck(clk), .q(\LUT[110][2] ) );
  dp_1 \LUT_reg[110][1]  ( .ip(n15227), .ck(clk), .q(\LUT[110][1] ) );
  dp_1 \LUT_reg[110][0]  ( .ip(n15226), .ck(clk), .q(\LUT[110][0] ) );
  dp_1 \LUT_reg[109][15]  ( .ip(n15225), .ck(clk), .q(\LUT[109][15] ) );
  dp_1 \LUT_reg[109][14]  ( .ip(n15224), .ck(clk), .q(\LUT[109][14] ) );
  dp_1 \LUT_reg[109][13]  ( .ip(n15223), .ck(clk), .q(\LUT[109][13] ) );
  dp_1 \LUT_reg[109][12]  ( .ip(n15222), .ck(clk), .q(\LUT[109][12] ) );
  dp_1 \LUT_reg[109][11]  ( .ip(n15221), .ck(clk), .q(\LUT[109][11] ) );
  dp_1 \LUT_reg[109][10]  ( .ip(n15220), .ck(clk), .q(\LUT[109][10] ) );
  dp_1 \LUT_reg[109][9]  ( .ip(n15219), .ck(clk), .q(\LUT[109][9] ) );
  dp_1 \LUT_reg[109][8]  ( .ip(n15218), .ck(clk), .q(\LUT[109][8] ) );
  dp_1 \LUT_reg[109][7]  ( .ip(n15217), .ck(clk), .q(\LUT[109][7] ) );
  dp_1 \LUT_reg[109][6]  ( .ip(n15216), .ck(clk), .q(\LUT[109][6] ) );
  dp_1 \LUT_reg[109][5]  ( .ip(n15215), .ck(clk), .q(\LUT[109][5] ) );
  dp_1 \LUT_reg[109][4]  ( .ip(n15214), .ck(clk), .q(\LUT[109][4] ) );
  dp_1 \LUT_reg[109][3]  ( .ip(n15213), .ck(clk), .q(\LUT[109][3] ) );
  dp_1 \LUT_reg[109][2]  ( .ip(n15212), .ck(clk), .q(\LUT[109][2] ) );
  dp_1 \LUT_reg[109][1]  ( .ip(n15211), .ck(clk), .q(\LUT[109][1] ) );
  dp_1 \LUT_reg[109][0]  ( .ip(n15210), .ck(clk), .q(\LUT[109][0] ) );
  dp_1 \LUT_reg[108][15]  ( .ip(n15209), .ck(clk), .q(\LUT[108][15] ) );
  dp_1 \LUT_reg[108][14]  ( .ip(n15208), .ck(clk), .q(\LUT[108][14] ) );
  dp_1 \LUT_reg[108][13]  ( .ip(n15207), .ck(clk), .q(\LUT[108][13] ) );
  dp_1 \LUT_reg[108][12]  ( .ip(n15206), .ck(clk), .q(\LUT[108][12] ) );
  dp_1 \LUT_reg[108][11]  ( .ip(n15205), .ck(clk), .q(\LUT[108][11] ) );
  dp_1 \LUT_reg[108][10]  ( .ip(n15204), .ck(clk), .q(\LUT[108][10] ) );
  dp_1 \LUT_reg[108][9]  ( .ip(n15203), .ck(clk), .q(\LUT[108][9] ) );
  dp_1 \LUT_reg[108][8]  ( .ip(n15202), .ck(clk), .q(\LUT[108][8] ) );
  dp_1 \LUT_reg[108][7]  ( .ip(n15201), .ck(clk), .q(\LUT[108][7] ) );
  dp_1 \LUT_reg[108][6]  ( .ip(n15200), .ck(clk), .q(\LUT[108][6] ) );
  dp_1 \LUT_reg[108][5]  ( .ip(n15199), .ck(clk), .q(\LUT[108][5] ) );
  dp_1 \LUT_reg[108][4]  ( .ip(n15198), .ck(clk), .q(\LUT[108][4] ) );
  dp_1 \LUT_reg[108][3]  ( .ip(n15197), .ck(clk), .q(\LUT[108][3] ) );
  dp_1 \LUT_reg[108][2]  ( .ip(n15196), .ck(clk), .q(\LUT[108][2] ) );
  dp_1 \LUT_reg[108][1]  ( .ip(n15195), .ck(clk), .q(\LUT[108][1] ) );
  dp_1 \LUT_reg[108][0]  ( .ip(n15194), .ck(clk), .q(\LUT[108][0] ) );
  dp_1 \LUT_reg[107][15]  ( .ip(n15193), .ck(clk), .q(\LUT[107][15] ) );
  dp_1 \LUT_reg[107][14]  ( .ip(n15192), .ck(clk), .q(\LUT[107][14] ) );
  dp_1 \LUT_reg[107][13]  ( .ip(n15191), .ck(clk), .q(\LUT[107][13] ) );
  dp_1 \LUT_reg[107][12]  ( .ip(n15190), .ck(clk), .q(\LUT[107][12] ) );
  dp_1 \LUT_reg[107][11]  ( .ip(n15189), .ck(clk), .q(\LUT[107][11] ) );
  dp_1 \LUT_reg[107][10]  ( .ip(n15188), .ck(clk), .q(\LUT[107][10] ) );
  dp_1 \LUT_reg[107][9]  ( .ip(n15187), .ck(clk), .q(\LUT[107][9] ) );
  dp_1 \LUT_reg[107][8]  ( .ip(n15186), .ck(clk), .q(\LUT[107][8] ) );
  dp_1 \LUT_reg[107][7]  ( .ip(n15185), .ck(clk), .q(\LUT[107][7] ) );
  dp_1 \LUT_reg[107][6]  ( .ip(n15184), .ck(clk), .q(\LUT[107][6] ) );
  dp_1 \LUT_reg[107][5]  ( .ip(n15183), .ck(clk), .q(\LUT[107][5] ) );
  dp_1 \LUT_reg[107][4]  ( .ip(n15182), .ck(clk), .q(\LUT[107][4] ) );
  dp_1 \LUT_reg[107][3]  ( .ip(n15181), .ck(clk), .q(\LUT[107][3] ) );
  dp_1 \LUT_reg[107][2]  ( .ip(n15180), .ck(clk), .q(\LUT[107][2] ) );
  dp_1 \LUT_reg[107][1]  ( .ip(n15179), .ck(clk), .q(\LUT[107][1] ) );
  dp_1 \LUT_reg[107][0]  ( .ip(n15178), .ck(clk), .q(\LUT[107][0] ) );
  dp_1 \LUT_reg[106][15]  ( .ip(n15177), .ck(clk), .q(\LUT[106][15] ) );
  dp_1 \LUT_reg[106][14]  ( .ip(n15176), .ck(clk), .q(\LUT[106][14] ) );
  dp_1 \LUT_reg[106][13]  ( .ip(n15175), .ck(clk), .q(\LUT[106][13] ) );
  dp_1 \LUT_reg[106][12]  ( .ip(n15174), .ck(clk), .q(\LUT[106][12] ) );
  dp_1 \LUT_reg[106][11]  ( .ip(n15173), .ck(clk), .q(\LUT[106][11] ) );
  dp_1 \LUT_reg[106][10]  ( .ip(n15172), .ck(clk), .q(\LUT[106][10] ) );
  dp_1 \LUT_reg[106][9]  ( .ip(n15171), .ck(clk), .q(\LUT[106][9] ) );
  dp_1 \LUT_reg[106][8]  ( .ip(n15170), .ck(clk), .q(\LUT[106][8] ) );
  dp_1 \LUT_reg[106][7]  ( .ip(n15169), .ck(clk), .q(\LUT[106][7] ) );
  dp_1 \LUT_reg[106][6]  ( .ip(n15168), .ck(clk), .q(\LUT[106][6] ) );
  dp_1 \LUT_reg[106][5]  ( .ip(n15167), .ck(clk), .q(\LUT[106][5] ) );
  dp_1 \LUT_reg[106][4]  ( .ip(n15166), .ck(clk), .q(\LUT[106][4] ) );
  dp_1 \LUT_reg[106][3]  ( .ip(n15165), .ck(clk), .q(\LUT[106][3] ) );
  dp_1 \LUT_reg[106][2]  ( .ip(n15164), .ck(clk), .q(\LUT[106][2] ) );
  dp_1 \LUT_reg[106][1]  ( .ip(n15163), .ck(clk), .q(\LUT[106][1] ) );
  dp_1 \LUT_reg[106][0]  ( .ip(n15162), .ck(clk), .q(\LUT[106][0] ) );
  dp_1 \LUT_reg[105][15]  ( .ip(n15161), .ck(clk), .q(\LUT[105][15] ) );
  dp_1 \LUT_reg[105][14]  ( .ip(n15160), .ck(clk), .q(\LUT[105][14] ) );
  dp_1 \LUT_reg[105][13]  ( .ip(n15159), .ck(clk), .q(\LUT[105][13] ) );
  dp_1 \LUT_reg[105][12]  ( .ip(n15158), .ck(clk), .q(\LUT[105][12] ) );
  dp_1 \LUT_reg[105][11]  ( .ip(n15157), .ck(clk), .q(\LUT[105][11] ) );
  dp_1 \LUT_reg[105][10]  ( .ip(n15156), .ck(clk), .q(\LUT[105][10] ) );
  dp_1 \LUT_reg[105][9]  ( .ip(n15155), .ck(clk), .q(\LUT[105][9] ) );
  dp_1 \LUT_reg[105][8]  ( .ip(n15154), .ck(clk), .q(\LUT[105][8] ) );
  dp_1 \LUT_reg[105][7]  ( .ip(n15153), .ck(clk), .q(\LUT[105][7] ) );
  dp_1 \LUT_reg[105][6]  ( .ip(n15152), .ck(clk), .q(\LUT[105][6] ) );
  dp_1 \LUT_reg[105][5]  ( .ip(n15151), .ck(clk), .q(\LUT[105][5] ) );
  dp_1 \LUT_reg[105][4]  ( .ip(n15150), .ck(clk), .q(\LUT[105][4] ) );
  dp_1 \LUT_reg[105][3]  ( .ip(n15149), .ck(clk), .q(\LUT[105][3] ) );
  dp_1 \LUT_reg[105][2]  ( .ip(n15148), .ck(clk), .q(\LUT[105][2] ) );
  dp_1 \LUT_reg[105][1]  ( .ip(n15147), .ck(clk), .q(\LUT[105][1] ) );
  dp_1 \LUT_reg[105][0]  ( .ip(n15146), .ck(clk), .q(\LUT[105][0] ) );
  dp_1 \LUT_reg[104][15]  ( .ip(n15145), .ck(clk), .q(\LUT[104][15] ) );
  dp_1 \LUT_reg[104][14]  ( .ip(n15144), .ck(clk), .q(\LUT[104][14] ) );
  dp_1 \LUT_reg[104][13]  ( .ip(n15143), .ck(clk), .q(\LUT[104][13] ) );
  dp_1 \LUT_reg[104][12]  ( .ip(n15142), .ck(clk), .q(\LUT[104][12] ) );
  dp_1 \LUT_reg[104][11]  ( .ip(n15141), .ck(clk), .q(\LUT[104][11] ) );
  dp_1 \LUT_reg[104][10]  ( .ip(n15140), .ck(clk), .q(\LUT[104][10] ) );
  dp_1 \LUT_reg[104][9]  ( .ip(n15139), .ck(clk), .q(\LUT[104][9] ) );
  dp_1 \LUT_reg[104][8]  ( .ip(n15138), .ck(clk), .q(\LUT[104][8] ) );
  dp_1 \LUT_reg[104][7]  ( .ip(n15137), .ck(clk), .q(\LUT[104][7] ) );
  dp_1 \LUT_reg[104][6]  ( .ip(n15136), .ck(clk), .q(\LUT[104][6] ) );
  dp_1 \LUT_reg[104][5]  ( .ip(n15135), .ck(clk), .q(\LUT[104][5] ) );
  dp_1 \LUT_reg[104][4]  ( .ip(n15134), .ck(clk), .q(\LUT[104][4] ) );
  dp_1 \LUT_reg[104][3]  ( .ip(n15133), .ck(clk), .q(\LUT[104][3] ) );
  dp_1 \LUT_reg[104][2]  ( .ip(n15132), .ck(clk), .q(\LUT[104][2] ) );
  dp_1 \LUT_reg[104][1]  ( .ip(n15131), .ck(clk), .q(\LUT[104][1] ) );
  dp_1 \LUT_reg[104][0]  ( .ip(n15130), .ck(clk), .q(\LUT[104][0] ) );
  dp_1 \LUT_reg[103][15]  ( .ip(n15129), .ck(clk), .q(\LUT[103][15] ) );
  dp_1 \LUT_reg[103][14]  ( .ip(n15128), .ck(clk), .q(\LUT[103][14] ) );
  dp_1 \LUT_reg[103][13]  ( .ip(n15127), .ck(clk), .q(\LUT[103][13] ) );
  dp_1 \LUT_reg[103][12]  ( .ip(n15126), .ck(clk), .q(\LUT[103][12] ) );
  dp_1 \LUT_reg[103][11]  ( .ip(n15125), .ck(clk), .q(\LUT[103][11] ) );
  dp_1 \LUT_reg[103][10]  ( .ip(n15124), .ck(clk), .q(\LUT[103][10] ) );
  dp_1 \LUT_reg[103][9]  ( .ip(n15123), .ck(clk), .q(\LUT[103][9] ) );
  dp_1 \LUT_reg[103][8]  ( .ip(n15122), .ck(clk), .q(\LUT[103][8] ) );
  dp_1 \LUT_reg[103][7]  ( .ip(n15121), .ck(clk), .q(\LUT[103][7] ) );
  dp_1 \LUT_reg[103][6]  ( .ip(n15120), .ck(clk), .q(\LUT[103][6] ) );
  dp_1 \LUT_reg[103][5]  ( .ip(n15119), .ck(clk), .q(\LUT[103][5] ) );
  dp_1 \LUT_reg[103][4]  ( .ip(n15118), .ck(clk), .q(\LUT[103][4] ) );
  dp_1 \LUT_reg[103][3]  ( .ip(n15117), .ck(clk), .q(\LUT[103][3] ) );
  dp_1 \LUT_reg[103][2]  ( .ip(n15116), .ck(clk), .q(\LUT[103][2] ) );
  dp_1 \LUT_reg[103][1]  ( .ip(n15115), .ck(clk), .q(\LUT[103][1] ) );
  dp_1 \LUT_reg[103][0]  ( .ip(n15114), .ck(clk), .q(\LUT[103][0] ) );
  dp_1 \LUT_reg[102][15]  ( .ip(n15113), .ck(clk), .q(\LUT[102][15] ) );
  dp_1 \LUT_reg[102][14]  ( .ip(n15112), .ck(clk), .q(\LUT[102][14] ) );
  dp_1 \LUT_reg[102][13]  ( .ip(n15111), .ck(clk), .q(\LUT[102][13] ) );
  dp_1 \LUT_reg[102][12]  ( .ip(n15110), .ck(clk), .q(\LUT[102][12] ) );
  dp_1 \LUT_reg[102][11]  ( .ip(n15109), .ck(clk), .q(\LUT[102][11] ) );
  dp_1 \LUT_reg[102][10]  ( .ip(n15108), .ck(clk), .q(\LUT[102][10] ) );
  dp_1 \LUT_reg[102][9]  ( .ip(n15107), .ck(clk), .q(\LUT[102][9] ) );
  dp_1 \LUT_reg[102][8]  ( .ip(n15106), .ck(clk), .q(\LUT[102][8] ) );
  dp_1 \LUT_reg[102][7]  ( .ip(n15105), .ck(clk), .q(\LUT[102][7] ) );
  dp_1 \LUT_reg[102][6]  ( .ip(n15104), .ck(clk), .q(\LUT[102][6] ) );
  dp_1 \LUT_reg[102][5]  ( .ip(n15103), .ck(clk), .q(\LUT[102][5] ) );
  dp_1 \LUT_reg[102][4]  ( .ip(n15102), .ck(clk), .q(\LUT[102][4] ) );
  dp_1 \LUT_reg[102][3]  ( .ip(n15101), .ck(clk), .q(\LUT[102][3] ) );
  dp_1 \LUT_reg[102][2]  ( .ip(n15100), .ck(clk), .q(\LUT[102][2] ) );
  dp_1 \LUT_reg[102][1]  ( .ip(n15099), .ck(clk), .q(\LUT[102][1] ) );
  dp_1 \LUT_reg[102][0]  ( .ip(n15098), .ck(clk), .q(\LUT[102][0] ) );
  dp_1 \LUT_reg[101][15]  ( .ip(n15097), .ck(clk), .q(\LUT[101][15] ) );
  dp_1 \LUT_reg[101][14]  ( .ip(n15096), .ck(clk), .q(\LUT[101][14] ) );
  dp_1 \LUT_reg[101][13]  ( .ip(n15095), .ck(clk), .q(\LUT[101][13] ) );
  dp_1 \LUT_reg[101][12]  ( .ip(n15094), .ck(clk), .q(\LUT[101][12] ) );
  dp_1 \LUT_reg[101][11]  ( .ip(n15093), .ck(clk), .q(\LUT[101][11] ) );
  dp_1 \LUT_reg[101][10]  ( .ip(n15092), .ck(clk), .q(\LUT[101][10] ) );
  dp_1 \LUT_reg[101][9]  ( .ip(n15091), .ck(clk), .q(\LUT[101][9] ) );
  dp_1 \LUT_reg[101][8]  ( .ip(n15090), .ck(clk), .q(\LUT[101][8] ) );
  dp_1 \LUT_reg[101][7]  ( .ip(n15089), .ck(clk), .q(\LUT[101][7] ) );
  dp_1 \LUT_reg[101][6]  ( .ip(n15088), .ck(clk), .q(\LUT[101][6] ) );
  dp_1 \LUT_reg[101][5]  ( .ip(n15087), .ck(clk), .q(\LUT[101][5] ) );
  dp_1 \LUT_reg[101][4]  ( .ip(n15086), .ck(clk), .q(\LUT[101][4] ) );
  dp_1 \LUT_reg[101][3]  ( .ip(n15085), .ck(clk), .q(\LUT[101][3] ) );
  dp_1 \LUT_reg[101][2]  ( .ip(n15084), .ck(clk), .q(\LUT[101][2] ) );
  dp_1 \LUT_reg[101][1]  ( .ip(n15083), .ck(clk), .q(\LUT[101][1] ) );
  dp_1 \LUT_reg[101][0]  ( .ip(n15082), .ck(clk), .q(\LUT[101][0] ) );
  dp_1 \LUT_reg[100][15]  ( .ip(n15081), .ck(clk), .q(\LUT[100][15] ) );
  dp_1 \LUT_reg[100][14]  ( .ip(n15080), .ck(clk), .q(\LUT[100][14] ) );
  dp_1 \LUT_reg[100][13]  ( .ip(n15079), .ck(clk), .q(\LUT[100][13] ) );
  dp_1 \LUT_reg[100][12]  ( .ip(n15078), .ck(clk), .q(\LUT[100][12] ) );
  dp_1 \LUT_reg[100][11]  ( .ip(n15077), .ck(clk), .q(\LUT[100][11] ) );
  dp_1 \LUT_reg[100][10]  ( .ip(n15076), .ck(clk), .q(\LUT[100][10] ) );
  dp_1 \LUT_reg[100][9]  ( .ip(n15075), .ck(clk), .q(\LUT[100][9] ) );
  dp_1 \LUT_reg[100][8]  ( .ip(n15074), .ck(clk), .q(\LUT[100][8] ) );
  dp_1 \LUT_reg[100][7]  ( .ip(n15073), .ck(clk), .q(\LUT[100][7] ) );
  dp_1 \LUT_reg[100][6]  ( .ip(n15072), .ck(clk), .q(\LUT[100][6] ) );
  dp_1 \LUT_reg[100][5]  ( .ip(n15071), .ck(clk), .q(\LUT[100][5] ) );
  dp_1 \LUT_reg[100][4]  ( .ip(n15070), .ck(clk), .q(\LUT[100][4] ) );
  dp_1 \LUT_reg[100][3]  ( .ip(n15069), .ck(clk), .q(\LUT[100][3] ) );
  dp_1 \LUT_reg[100][2]  ( .ip(n15068), .ck(clk), .q(\LUT[100][2] ) );
  dp_1 \LUT_reg[100][1]  ( .ip(n15067), .ck(clk), .q(\LUT[100][1] ) );
  dp_1 \LUT_reg[100][0]  ( .ip(n15066), .ck(clk), .q(\LUT[100][0] ) );
  dp_1 \LUT_reg[99][15]  ( .ip(n15065), .ck(clk), .q(\LUT[99][15] ) );
  dp_1 \LUT_reg[99][14]  ( .ip(n15064), .ck(clk), .q(\LUT[99][14] ) );
  dp_1 \LUT_reg[99][13]  ( .ip(n15063), .ck(clk), .q(\LUT[99][13] ) );
  dp_1 \LUT_reg[99][12]  ( .ip(n15062), .ck(clk), .q(\LUT[99][12] ) );
  dp_1 \LUT_reg[99][11]  ( .ip(n15061), .ck(clk), .q(\LUT[99][11] ) );
  dp_1 \LUT_reg[99][10]  ( .ip(n15060), .ck(clk), .q(\LUT[99][10] ) );
  dp_1 \LUT_reg[99][9]  ( .ip(n15059), .ck(clk), .q(\LUT[99][9] ) );
  dp_1 \LUT_reg[99][8]  ( .ip(n15058), .ck(clk), .q(\LUT[99][8] ) );
  dp_1 \LUT_reg[99][7]  ( .ip(n15057), .ck(clk), .q(\LUT[99][7] ) );
  dp_1 \LUT_reg[99][6]  ( .ip(n15056), .ck(clk), .q(\LUT[99][6] ) );
  dp_1 \LUT_reg[99][5]  ( .ip(n15055), .ck(clk), .q(\LUT[99][5] ) );
  dp_1 \LUT_reg[99][4]  ( .ip(n15054), .ck(clk), .q(\LUT[99][4] ) );
  dp_1 \LUT_reg[99][3]  ( .ip(n15053), .ck(clk), .q(\LUT[99][3] ) );
  dp_1 \LUT_reg[99][2]  ( .ip(n15052), .ck(clk), .q(\LUT[99][2] ) );
  dp_1 \LUT_reg[99][1]  ( .ip(n15051), .ck(clk), .q(\LUT[99][1] ) );
  dp_1 \LUT_reg[99][0]  ( .ip(n15050), .ck(clk), .q(\LUT[99][0] ) );
  dp_1 \LUT_reg[98][15]  ( .ip(n15049), .ck(clk), .q(\LUT[98][15] ) );
  dp_1 \LUT_reg[98][14]  ( .ip(n15048), .ck(clk), .q(\LUT[98][14] ) );
  dp_1 \LUT_reg[98][13]  ( .ip(n15047), .ck(clk), .q(\LUT[98][13] ) );
  dp_1 \LUT_reg[98][12]  ( .ip(n15046), .ck(clk), .q(\LUT[98][12] ) );
  dp_1 \LUT_reg[98][11]  ( .ip(n15045), .ck(clk), .q(\LUT[98][11] ) );
  dp_1 \LUT_reg[98][10]  ( .ip(n15044), .ck(clk), .q(\LUT[98][10] ) );
  dp_1 \LUT_reg[98][9]  ( .ip(n15043), .ck(clk), .q(\LUT[98][9] ) );
  dp_1 \LUT_reg[98][8]  ( .ip(n15042), .ck(clk), .q(\LUT[98][8] ) );
  dp_1 \LUT_reg[98][7]  ( .ip(n15041), .ck(clk), .q(\LUT[98][7] ) );
  dp_1 \LUT_reg[98][6]  ( .ip(n15040), .ck(clk), .q(\LUT[98][6] ) );
  dp_1 \LUT_reg[98][5]  ( .ip(n15039), .ck(clk), .q(\LUT[98][5] ) );
  dp_1 \LUT_reg[98][4]  ( .ip(n15038), .ck(clk), .q(\LUT[98][4] ) );
  dp_1 \LUT_reg[98][3]  ( .ip(n15037), .ck(clk), .q(\LUT[98][3] ) );
  dp_1 \LUT_reg[98][2]  ( .ip(n15036), .ck(clk), .q(\LUT[98][2] ) );
  dp_1 \LUT_reg[98][1]  ( .ip(n15035), .ck(clk), .q(\LUT[98][1] ) );
  dp_1 \LUT_reg[98][0]  ( .ip(n15034), .ck(clk), .q(\LUT[98][0] ) );
  dp_1 \LUT_reg[97][15]  ( .ip(n15033), .ck(clk), .q(\LUT[97][15] ) );
  dp_1 \LUT_reg[97][14]  ( .ip(n15032), .ck(clk), .q(\LUT[97][14] ) );
  dp_1 \LUT_reg[97][13]  ( .ip(n15031), .ck(clk), .q(\LUT[97][13] ) );
  dp_1 \LUT_reg[97][12]  ( .ip(n15030), .ck(clk), .q(\LUT[97][12] ) );
  dp_1 \LUT_reg[97][11]  ( .ip(n15029), .ck(clk), .q(\LUT[97][11] ) );
  dp_1 \LUT_reg[97][10]  ( .ip(n15028), .ck(clk), .q(\LUT[97][10] ) );
  dp_1 \LUT_reg[97][9]  ( .ip(n15027), .ck(clk), .q(\LUT[97][9] ) );
  dp_1 \LUT_reg[97][8]  ( .ip(n15026), .ck(clk), .q(\LUT[97][8] ) );
  dp_1 \LUT_reg[97][7]  ( .ip(n15025), .ck(clk), .q(\LUT[97][7] ) );
  dp_1 \LUT_reg[97][6]  ( .ip(n15024), .ck(clk), .q(\LUT[97][6] ) );
  dp_1 \LUT_reg[97][5]  ( .ip(n15023), .ck(clk), .q(\LUT[97][5] ) );
  dp_1 \LUT_reg[97][4]  ( .ip(n15022), .ck(clk), .q(\LUT[97][4] ) );
  dp_1 \LUT_reg[97][3]  ( .ip(n15021), .ck(clk), .q(\LUT[97][3] ) );
  dp_1 \LUT_reg[97][2]  ( .ip(n15020), .ck(clk), .q(\LUT[97][2] ) );
  dp_1 \LUT_reg[97][1]  ( .ip(n15019), .ck(clk), .q(\LUT[97][1] ) );
  dp_1 \LUT_reg[97][0]  ( .ip(n15018), .ck(clk), .q(\LUT[97][0] ) );
  dp_1 \LUT_reg[96][15]  ( .ip(n15017), .ck(clk), .q(\LUT[96][15] ) );
  dp_1 \LUT_reg[96][14]  ( .ip(n15016), .ck(clk), .q(\LUT[96][14] ) );
  dp_1 \LUT_reg[96][13]  ( .ip(n15015), .ck(clk), .q(\LUT[96][13] ) );
  dp_1 \LUT_reg[96][12]  ( .ip(n15014), .ck(clk), .q(\LUT[96][12] ) );
  dp_1 \LUT_reg[96][11]  ( .ip(n15013), .ck(clk), .q(\LUT[96][11] ) );
  dp_1 \LUT_reg[96][10]  ( .ip(n15012), .ck(clk), .q(\LUT[96][10] ) );
  dp_1 \LUT_reg[96][9]  ( .ip(n15011), .ck(clk), .q(\LUT[96][9] ) );
  dp_1 \LUT_reg[96][8]  ( .ip(n15010), .ck(clk), .q(\LUT[96][8] ) );
  dp_1 \LUT_reg[96][7]  ( .ip(n15009), .ck(clk), .q(\LUT[96][7] ) );
  dp_1 \LUT_reg[96][6]  ( .ip(n15008), .ck(clk), .q(\LUT[96][6] ) );
  dp_1 \LUT_reg[96][5]  ( .ip(n15007), .ck(clk), .q(\LUT[96][5] ) );
  dp_1 \LUT_reg[96][4]  ( .ip(n15006), .ck(clk), .q(\LUT[96][4] ) );
  dp_1 \LUT_reg[96][3]  ( .ip(n15005), .ck(clk), .q(\LUT[96][3] ) );
  dp_1 \LUT_reg[96][2]  ( .ip(n15004), .ck(clk), .q(\LUT[96][2] ) );
  dp_1 \LUT_reg[96][1]  ( .ip(n15003), .ck(clk), .q(\LUT[96][1] ) );
  dp_1 \LUT_reg[96][0]  ( .ip(n15002), .ck(clk), .q(\LUT[96][0] ) );
  dp_1 \LUT_reg[95][15]  ( .ip(n15001), .ck(clk), .q(\LUT[95][15] ) );
  dp_1 \LUT_reg[95][14]  ( .ip(n15000), .ck(clk), .q(\LUT[95][14] ) );
  dp_1 \LUT_reg[95][13]  ( .ip(n14999), .ck(clk), .q(\LUT[95][13] ) );
  dp_1 \LUT_reg[95][12]  ( .ip(n14998), .ck(clk), .q(\LUT[95][12] ) );
  dp_1 \LUT_reg[95][11]  ( .ip(n14997), .ck(clk), .q(\LUT[95][11] ) );
  dp_1 \LUT_reg[95][10]  ( .ip(n14996), .ck(clk), .q(\LUT[95][10] ) );
  dp_1 \LUT_reg[95][9]  ( .ip(n14995), .ck(clk), .q(\LUT[95][9] ) );
  dp_1 \LUT_reg[95][8]  ( .ip(n14994), .ck(clk), .q(\LUT[95][8] ) );
  dp_1 \LUT_reg[95][7]  ( .ip(n14993), .ck(clk), .q(\LUT[95][7] ) );
  dp_1 \LUT_reg[95][6]  ( .ip(n14992), .ck(clk), .q(\LUT[95][6] ) );
  dp_1 \LUT_reg[95][5]  ( .ip(n14991), .ck(clk), .q(\LUT[95][5] ) );
  dp_1 \LUT_reg[95][4]  ( .ip(n14990), .ck(clk), .q(\LUT[95][4] ) );
  dp_1 \LUT_reg[95][3]  ( .ip(n14989), .ck(clk), .q(\LUT[95][3] ) );
  dp_1 \LUT_reg[95][2]  ( .ip(n14988), .ck(clk), .q(\LUT[95][2] ) );
  dp_1 \LUT_reg[95][1]  ( .ip(n14987), .ck(clk), .q(\LUT[95][1] ) );
  dp_1 \LUT_reg[95][0]  ( .ip(n14986), .ck(clk), .q(\LUT[95][0] ) );
  dp_1 \LUT_reg[94][15]  ( .ip(n14985), .ck(clk), .q(\LUT[94][15] ) );
  dp_1 \LUT_reg[94][14]  ( .ip(n14984), .ck(clk), .q(\LUT[94][14] ) );
  dp_1 \LUT_reg[94][13]  ( .ip(n14983), .ck(clk), .q(\LUT[94][13] ) );
  dp_1 \LUT_reg[94][12]  ( .ip(n14982), .ck(clk), .q(\LUT[94][12] ) );
  dp_1 \LUT_reg[94][11]  ( .ip(n14981), .ck(clk), .q(\LUT[94][11] ) );
  dp_1 \LUT_reg[94][10]  ( .ip(n14980), .ck(clk), .q(\LUT[94][10] ) );
  dp_1 \LUT_reg[94][9]  ( .ip(n14979), .ck(clk), .q(\LUT[94][9] ) );
  dp_1 \LUT_reg[94][8]  ( .ip(n14978), .ck(clk), .q(\LUT[94][8] ) );
  dp_1 \LUT_reg[94][7]  ( .ip(n14977), .ck(clk), .q(\LUT[94][7] ) );
  dp_1 \LUT_reg[94][6]  ( .ip(n14976), .ck(clk), .q(\LUT[94][6] ) );
  dp_1 \LUT_reg[94][5]  ( .ip(n14975), .ck(clk), .q(\LUT[94][5] ) );
  dp_1 \LUT_reg[94][4]  ( .ip(n14974), .ck(clk), .q(\LUT[94][4] ) );
  dp_1 \LUT_reg[94][3]  ( .ip(n14973), .ck(clk), .q(\LUT[94][3] ) );
  dp_1 \LUT_reg[94][2]  ( .ip(n14972), .ck(clk), .q(\LUT[94][2] ) );
  dp_1 \LUT_reg[94][1]  ( .ip(n14971), .ck(clk), .q(\LUT[94][1] ) );
  dp_1 \LUT_reg[94][0]  ( .ip(n14970), .ck(clk), .q(\LUT[94][0] ) );
  dp_1 \LUT_reg[93][15]  ( .ip(n14969), .ck(clk), .q(\LUT[93][15] ) );
  dp_1 \LUT_reg[93][14]  ( .ip(n14968), .ck(clk), .q(\LUT[93][14] ) );
  dp_1 \LUT_reg[93][13]  ( .ip(n14967), .ck(clk), .q(\LUT[93][13] ) );
  dp_1 \LUT_reg[93][12]  ( .ip(n14966), .ck(clk), .q(\LUT[93][12] ) );
  dp_1 \LUT_reg[93][11]  ( .ip(n14965), .ck(clk), .q(\LUT[93][11] ) );
  dp_1 \LUT_reg[93][10]  ( .ip(n14964), .ck(clk), .q(\LUT[93][10] ) );
  dp_1 \LUT_reg[93][9]  ( .ip(n14963), .ck(clk), .q(\LUT[93][9] ) );
  dp_1 \LUT_reg[93][8]  ( .ip(n14962), .ck(clk), .q(\LUT[93][8] ) );
  dp_1 \LUT_reg[93][7]  ( .ip(n14961), .ck(clk), .q(\LUT[93][7] ) );
  dp_1 \LUT_reg[93][6]  ( .ip(n14960), .ck(clk), .q(\LUT[93][6] ) );
  dp_1 \LUT_reg[93][5]  ( .ip(n14959), .ck(clk), .q(\LUT[93][5] ) );
  dp_1 \LUT_reg[93][4]  ( .ip(n14958), .ck(clk), .q(\LUT[93][4] ) );
  dp_1 \LUT_reg[93][3]  ( .ip(n14957), .ck(clk), .q(\LUT[93][3] ) );
  dp_1 \LUT_reg[93][2]  ( .ip(n14956), .ck(clk), .q(\LUT[93][2] ) );
  dp_1 \LUT_reg[93][1]  ( .ip(n14955), .ck(clk), .q(\LUT[93][1] ) );
  dp_1 \LUT_reg[93][0]  ( .ip(n14954), .ck(clk), .q(\LUT[93][0] ) );
  dp_1 \LUT_reg[92][15]  ( .ip(n14953), .ck(clk), .q(\LUT[92][15] ) );
  dp_1 \LUT_reg[92][14]  ( .ip(n14952), .ck(clk), .q(\LUT[92][14] ) );
  dp_1 \LUT_reg[92][13]  ( .ip(n14951), .ck(clk), .q(\LUT[92][13] ) );
  dp_1 \LUT_reg[92][12]  ( .ip(n14950), .ck(clk), .q(\LUT[92][12] ) );
  dp_1 \LUT_reg[92][11]  ( .ip(n14949), .ck(clk), .q(\LUT[92][11] ) );
  dp_1 \LUT_reg[92][10]  ( .ip(n14948), .ck(clk), .q(\LUT[92][10] ) );
  dp_1 \LUT_reg[92][9]  ( .ip(n14947), .ck(clk), .q(\LUT[92][9] ) );
  dp_1 \LUT_reg[92][8]  ( .ip(n14946), .ck(clk), .q(\LUT[92][8] ) );
  dp_1 \LUT_reg[92][7]  ( .ip(n14945), .ck(clk), .q(\LUT[92][7] ) );
  dp_1 \LUT_reg[92][6]  ( .ip(n14944), .ck(clk), .q(\LUT[92][6] ) );
  dp_1 \LUT_reg[92][5]  ( .ip(n14943), .ck(clk), .q(\LUT[92][5] ) );
  dp_1 \LUT_reg[92][4]  ( .ip(n14942), .ck(clk), .q(\LUT[92][4] ) );
  dp_1 \LUT_reg[92][3]  ( .ip(n14941), .ck(clk), .q(\LUT[92][3] ) );
  dp_1 \LUT_reg[92][2]  ( .ip(n14940), .ck(clk), .q(\LUT[92][2] ) );
  dp_1 \LUT_reg[92][1]  ( .ip(n14939), .ck(clk), .q(\LUT[92][1] ) );
  dp_1 \LUT_reg[92][0]  ( .ip(n14938), .ck(clk), .q(\LUT[92][0] ) );
  dp_1 \LUT_reg[91][15]  ( .ip(n14937), .ck(clk), .q(\LUT[91][15] ) );
  dp_1 \LUT_reg[91][14]  ( .ip(n14936), .ck(clk), .q(\LUT[91][14] ) );
  dp_1 \LUT_reg[91][13]  ( .ip(n14935), .ck(clk), .q(\LUT[91][13] ) );
  dp_1 \LUT_reg[91][12]  ( .ip(n14934), .ck(clk), .q(\LUT[91][12] ) );
  dp_1 \LUT_reg[91][11]  ( .ip(n14933), .ck(clk), .q(\LUT[91][11] ) );
  dp_1 \LUT_reg[91][10]  ( .ip(n14932), .ck(clk), .q(\LUT[91][10] ) );
  dp_1 \LUT_reg[91][9]  ( .ip(n14931), .ck(clk), .q(\LUT[91][9] ) );
  dp_1 \LUT_reg[91][8]  ( .ip(n14930), .ck(clk), .q(\LUT[91][8] ) );
  dp_1 \LUT_reg[91][7]  ( .ip(n14929), .ck(clk), .q(\LUT[91][7] ) );
  dp_1 \LUT_reg[91][6]  ( .ip(n14928), .ck(clk), .q(\LUT[91][6] ) );
  dp_1 \LUT_reg[91][5]  ( .ip(n14927), .ck(clk), .q(\LUT[91][5] ) );
  dp_1 \LUT_reg[91][4]  ( .ip(n14926), .ck(clk), .q(\LUT[91][4] ) );
  dp_1 \LUT_reg[91][3]  ( .ip(n14925), .ck(clk), .q(\LUT[91][3] ) );
  dp_1 \LUT_reg[91][2]  ( .ip(n14924), .ck(clk), .q(\LUT[91][2] ) );
  dp_1 \LUT_reg[91][1]  ( .ip(n14923), .ck(clk), .q(\LUT[91][1] ) );
  dp_1 \LUT_reg[91][0]  ( .ip(n14922), .ck(clk), .q(\LUT[91][0] ) );
  dp_1 \LUT_reg[90][15]  ( .ip(n14921), .ck(clk), .q(\LUT[90][15] ) );
  dp_1 \LUT_reg[90][14]  ( .ip(n14920), .ck(clk), .q(\LUT[90][14] ) );
  dp_1 \LUT_reg[90][13]  ( .ip(n14919), .ck(clk), .q(\LUT[90][13] ) );
  dp_1 \LUT_reg[90][12]  ( .ip(n14918), .ck(clk), .q(\LUT[90][12] ) );
  dp_1 \LUT_reg[90][11]  ( .ip(n14917), .ck(clk), .q(\LUT[90][11] ) );
  dp_1 \LUT_reg[90][10]  ( .ip(n14916), .ck(clk), .q(\LUT[90][10] ) );
  dp_1 \LUT_reg[90][9]  ( .ip(n14915), .ck(clk), .q(\LUT[90][9] ) );
  dp_1 \LUT_reg[90][8]  ( .ip(n14914), .ck(clk), .q(\LUT[90][8] ) );
  dp_1 \LUT_reg[90][7]  ( .ip(n14913), .ck(clk), .q(\LUT[90][7] ) );
  dp_1 \LUT_reg[90][6]  ( .ip(n14912), .ck(clk), .q(\LUT[90][6] ) );
  dp_1 \LUT_reg[90][5]  ( .ip(n14911), .ck(clk), .q(\LUT[90][5] ) );
  dp_1 \LUT_reg[90][4]  ( .ip(n14910), .ck(clk), .q(\LUT[90][4] ) );
  dp_1 \LUT_reg[90][3]  ( .ip(n14909), .ck(clk), .q(\LUT[90][3] ) );
  dp_1 \LUT_reg[90][2]  ( .ip(n14908), .ck(clk), .q(\LUT[90][2] ) );
  dp_1 \LUT_reg[90][1]  ( .ip(n14907), .ck(clk), .q(\LUT[90][1] ) );
  dp_1 \LUT_reg[90][0]  ( .ip(n14906), .ck(clk), .q(\LUT[90][0] ) );
  dp_1 \LUT_reg[89][15]  ( .ip(n14905), .ck(clk), .q(\LUT[89][15] ) );
  dp_1 \LUT_reg[89][14]  ( .ip(n14904), .ck(clk), .q(\LUT[89][14] ) );
  dp_1 \LUT_reg[89][13]  ( .ip(n14903), .ck(clk), .q(\LUT[89][13] ) );
  dp_1 \LUT_reg[89][12]  ( .ip(n14902), .ck(clk), .q(\LUT[89][12] ) );
  dp_1 \LUT_reg[89][11]  ( .ip(n14901), .ck(clk), .q(\LUT[89][11] ) );
  dp_1 \LUT_reg[89][10]  ( .ip(n14900), .ck(clk), .q(\LUT[89][10] ) );
  dp_1 \LUT_reg[89][9]  ( .ip(n14899), .ck(clk), .q(\LUT[89][9] ) );
  dp_1 \LUT_reg[89][8]  ( .ip(n14898), .ck(clk), .q(\LUT[89][8] ) );
  dp_1 \LUT_reg[89][7]  ( .ip(n14897), .ck(clk), .q(\LUT[89][7] ) );
  dp_1 \LUT_reg[89][6]  ( .ip(n14896), .ck(clk), .q(\LUT[89][6] ) );
  dp_1 \LUT_reg[89][5]  ( .ip(n14895), .ck(clk), .q(\LUT[89][5] ) );
  dp_1 \LUT_reg[89][4]  ( .ip(n14894), .ck(clk), .q(\LUT[89][4] ) );
  dp_1 \LUT_reg[89][3]  ( .ip(n14893), .ck(clk), .q(\LUT[89][3] ) );
  dp_1 \LUT_reg[89][2]  ( .ip(n14892), .ck(clk), .q(\LUT[89][2] ) );
  dp_1 \LUT_reg[89][1]  ( .ip(n14891), .ck(clk), .q(\LUT[89][1] ) );
  dp_1 \LUT_reg[89][0]  ( .ip(n14890), .ck(clk), .q(\LUT[89][0] ) );
  dp_1 \LUT_reg[88][15]  ( .ip(n14889), .ck(clk), .q(\LUT[88][15] ) );
  dp_1 \LUT_reg[88][14]  ( .ip(n14888), .ck(clk), .q(\LUT[88][14] ) );
  dp_1 \LUT_reg[88][13]  ( .ip(n14887), .ck(clk), .q(\LUT[88][13] ) );
  dp_1 \LUT_reg[88][12]  ( .ip(n14886), .ck(clk), .q(\LUT[88][12] ) );
  dp_1 \LUT_reg[88][11]  ( .ip(n14885), .ck(clk), .q(\LUT[88][11] ) );
  dp_1 \LUT_reg[88][10]  ( .ip(n14884), .ck(clk), .q(\LUT[88][10] ) );
  dp_1 \LUT_reg[88][9]  ( .ip(n14883), .ck(clk), .q(\LUT[88][9] ) );
  dp_1 \LUT_reg[88][8]  ( .ip(n14882), .ck(clk), .q(\LUT[88][8] ) );
  dp_1 \LUT_reg[88][7]  ( .ip(n14881), .ck(clk), .q(\LUT[88][7] ) );
  dp_1 \LUT_reg[88][6]  ( .ip(n14880), .ck(clk), .q(\LUT[88][6] ) );
  dp_1 \LUT_reg[88][5]  ( .ip(n14879), .ck(clk), .q(\LUT[88][5] ) );
  dp_1 \LUT_reg[88][4]  ( .ip(n14878), .ck(clk), .q(\LUT[88][4] ) );
  dp_1 \LUT_reg[88][3]  ( .ip(n14877), .ck(clk), .q(\LUT[88][3] ) );
  dp_1 \LUT_reg[88][2]  ( .ip(n14876), .ck(clk), .q(\LUT[88][2] ) );
  dp_1 \LUT_reg[88][1]  ( .ip(n14875), .ck(clk), .q(\LUT[88][1] ) );
  dp_1 \LUT_reg[88][0]  ( .ip(n14874), .ck(clk), .q(\LUT[88][0] ) );
  dp_1 \LUT_reg[87][15]  ( .ip(n14873), .ck(clk), .q(\LUT[87][15] ) );
  dp_1 \LUT_reg[87][14]  ( .ip(n14872), .ck(clk), .q(\LUT[87][14] ) );
  dp_1 \LUT_reg[87][13]  ( .ip(n14871), .ck(clk), .q(\LUT[87][13] ) );
  dp_1 \LUT_reg[87][12]  ( .ip(n14870), .ck(clk), .q(\LUT[87][12] ) );
  dp_1 \LUT_reg[87][11]  ( .ip(n14869), .ck(clk), .q(\LUT[87][11] ) );
  dp_1 \LUT_reg[87][10]  ( .ip(n14868), .ck(clk), .q(\LUT[87][10] ) );
  dp_1 \LUT_reg[87][9]  ( .ip(n14867), .ck(clk), .q(\LUT[87][9] ) );
  dp_1 \LUT_reg[87][8]  ( .ip(n14866), .ck(clk), .q(\LUT[87][8] ) );
  dp_1 \LUT_reg[87][7]  ( .ip(n14865), .ck(clk), .q(\LUT[87][7] ) );
  dp_1 \LUT_reg[87][6]  ( .ip(n14864), .ck(clk), .q(\LUT[87][6] ) );
  dp_1 \LUT_reg[87][5]  ( .ip(n14863), .ck(clk), .q(\LUT[87][5] ) );
  dp_1 \LUT_reg[87][4]  ( .ip(n14862), .ck(clk), .q(\LUT[87][4] ) );
  dp_1 \LUT_reg[87][3]  ( .ip(n14861), .ck(clk), .q(\LUT[87][3] ) );
  dp_1 \LUT_reg[87][2]  ( .ip(n14860), .ck(clk), .q(\LUT[87][2] ) );
  dp_1 \LUT_reg[87][1]  ( .ip(n14859), .ck(clk), .q(\LUT[87][1] ) );
  dp_1 \LUT_reg[87][0]  ( .ip(n14858), .ck(clk), .q(\LUT[87][0] ) );
  dp_1 \LUT_reg[86][15]  ( .ip(n14857), .ck(clk), .q(\LUT[86][15] ) );
  dp_1 \LUT_reg[86][14]  ( .ip(n14856), .ck(clk), .q(\LUT[86][14] ) );
  dp_1 \LUT_reg[86][13]  ( .ip(n14855), .ck(clk), .q(\LUT[86][13] ) );
  dp_1 \LUT_reg[86][12]  ( .ip(n14854), .ck(clk), .q(\LUT[86][12] ) );
  dp_1 \LUT_reg[86][11]  ( .ip(n14853), .ck(clk), .q(\LUT[86][11] ) );
  dp_1 \LUT_reg[86][10]  ( .ip(n14852), .ck(clk), .q(\LUT[86][10] ) );
  dp_1 \LUT_reg[86][9]  ( .ip(n14851), .ck(clk), .q(\LUT[86][9] ) );
  dp_1 \LUT_reg[86][8]  ( .ip(n14850), .ck(clk), .q(\LUT[86][8] ) );
  dp_1 \LUT_reg[86][7]  ( .ip(n14849), .ck(clk), .q(\LUT[86][7] ) );
  dp_1 \LUT_reg[86][6]  ( .ip(n14848), .ck(clk), .q(\LUT[86][6] ) );
  dp_1 \LUT_reg[86][5]  ( .ip(n14847), .ck(clk), .q(\LUT[86][5] ) );
  dp_1 \LUT_reg[86][4]  ( .ip(n14846), .ck(clk), .q(\LUT[86][4] ) );
  dp_1 \LUT_reg[86][3]  ( .ip(n14845), .ck(clk), .q(\LUT[86][3] ) );
  dp_1 \LUT_reg[86][2]  ( .ip(n14844), .ck(clk), .q(\LUT[86][2] ) );
  dp_1 \LUT_reg[86][1]  ( .ip(n14843), .ck(clk), .q(\LUT[86][1] ) );
  dp_1 \LUT_reg[86][0]  ( .ip(n14842), .ck(clk), .q(\LUT[86][0] ) );
  dp_1 \LUT_reg[85][15]  ( .ip(n14841), .ck(clk), .q(\LUT[85][15] ) );
  dp_1 \LUT_reg[85][14]  ( .ip(n14840), .ck(clk), .q(\LUT[85][14] ) );
  dp_1 \LUT_reg[85][13]  ( .ip(n14839), .ck(clk), .q(\LUT[85][13] ) );
  dp_1 \LUT_reg[85][12]  ( .ip(n14838), .ck(clk), .q(\LUT[85][12] ) );
  dp_1 \LUT_reg[85][11]  ( .ip(n14837), .ck(clk), .q(\LUT[85][11] ) );
  dp_1 \LUT_reg[85][10]  ( .ip(n14836), .ck(clk), .q(\LUT[85][10] ) );
  dp_1 \LUT_reg[85][9]  ( .ip(n14835), .ck(clk), .q(\LUT[85][9] ) );
  dp_1 \LUT_reg[85][8]  ( .ip(n14834), .ck(clk), .q(\LUT[85][8] ) );
  dp_1 \LUT_reg[85][7]  ( .ip(n14833), .ck(clk), .q(\LUT[85][7] ) );
  dp_1 \LUT_reg[85][6]  ( .ip(n14832), .ck(clk), .q(\LUT[85][6] ) );
  dp_1 \LUT_reg[85][5]  ( .ip(n14831), .ck(clk), .q(\LUT[85][5] ) );
  dp_1 \LUT_reg[85][4]  ( .ip(n14830), .ck(clk), .q(\LUT[85][4] ) );
  dp_1 \LUT_reg[85][3]  ( .ip(n14829), .ck(clk), .q(\LUT[85][3] ) );
  dp_1 \LUT_reg[85][2]  ( .ip(n14828), .ck(clk), .q(\LUT[85][2] ) );
  dp_1 \LUT_reg[85][1]  ( .ip(n14827), .ck(clk), .q(\LUT[85][1] ) );
  dp_1 \LUT_reg[85][0]  ( .ip(n14826), .ck(clk), .q(\LUT[85][0] ) );
  dp_1 \LUT_reg[84][15]  ( .ip(n14825), .ck(clk), .q(\LUT[84][15] ) );
  dp_1 \LUT_reg[84][14]  ( .ip(n14824), .ck(clk), .q(\LUT[84][14] ) );
  dp_1 \LUT_reg[84][13]  ( .ip(n14823), .ck(clk), .q(\LUT[84][13] ) );
  dp_1 \LUT_reg[84][12]  ( .ip(n14822), .ck(clk), .q(\LUT[84][12] ) );
  dp_1 \LUT_reg[84][11]  ( .ip(n14821), .ck(clk), .q(\LUT[84][11] ) );
  dp_1 \LUT_reg[84][10]  ( .ip(n14820), .ck(clk), .q(\LUT[84][10] ) );
  dp_1 \LUT_reg[84][9]  ( .ip(n14819), .ck(clk), .q(\LUT[84][9] ) );
  dp_1 \LUT_reg[84][8]  ( .ip(n14818), .ck(clk), .q(\LUT[84][8] ) );
  dp_1 \LUT_reg[84][7]  ( .ip(n14817), .ck(clk), .q(\LUT[84][7] ) );
  dp_1 \LUT_reg[84][6]  ( .ip(n14816), .ck(clk), .q(\LUT[84][6] ) );
  dp_1 \LUT_reg[84][5]  ( .ip(n14815), .ck(clk), .q(\LUT[84][5] ) );
  dp_1 \LUT_reg[84][4]  ( .ip(n14814), .ck(clk), .q(\LUT[84][4] ) );
  dp_1 \LUT_reg[84][3]  ( .ip(n14813), .ck(clk), .q(\LUT[84][3] ) );
  dp_1 \LUT_reg[84][2]  ( .ip(n14812), .ck(clk), .q(\LUT[84][2] ) );
  dp_1 \LUT_reg[84][1]  ( .ip(n14811), .ck(clk), .q(\LUT[84][1] ) );
  dp_1 \LUT_reg[84][0]  ( .ip(n14810), .ck(clk), .q(\LUT[84][0] ) );
  dp_1 \LUT_reg[83][15]  ( .ip(n14809), .ck(clk), .q(\LUT[83][15] ) );
  dp_1 \LUT_reg[83][14]  ( .ip(n14808), .ck(clk), .q(\LUT[83][14] ) );
  dp_1 \LUT_reg[83][13]  ( .ip(n14807), .ck(clk), .q(\LUT[83][13] ) );
  dp_1 \LUT_reg[83][12]  ( .ip(n14806), .ck(clk), .q(\LUT[83][12] ) );
  dp_1 \LUT_reg[83][11]  ( .ip(n14805), .ck(clk), .q(\LUT[83][11] ) );
  dp_1 \LUT_reg[83][10]  ( .ip(n14804), .ck(clk), .q(\LUT[83][10] ) );
  dp_1 \LUT_reg[83][9]  ( .ip(n14803), .ck(clk), .q(\LUT[83][9] ) );
  dp_1 \LUT_reg[83][8]  ( .ip(n14802), .ck(clk), .q(\LUT[83][8] ) );
  dp_1 \LUT_reg[83][7]  ( .ip(n14801), .ck(clk), .q(\LUT[83][7] ) );
  dp_1 \LUT_reg[83][6]  ( .ip(n14800), .ck(clk), .q(\LUT[83][6] ) );
  dp_1 \LUT_reg[83][5]  ( .ip(n14799), .ck(clk), .q(\LUT[83][5] ) );
  dp_1 \LUT_reg[83][4]  ( .ip(n14798), .ck(clk), .q(\LUT[83][4] ) );
  dp_1 \LUT_reg[83][3]  ( .ip(n14797), .ck(clk), .q(\LUT[83][3] ) );
  dp_1 \LUT_reg[83][2]  ( .ip(n14796), .ck(clk), .q(\LUT[83][2] ) );
  dp_1 \LUT_reg[83][1]  ( .ip(n14795), .ck(clk), .q(\LUT[83][1] ) );
  dp_1 \LUT_reg[83][0]  ( .ip(n14794), .ck(clk), .q(\LUT[83][0] ) );
  dp_1 \LUT_reg[82][15]  ( .ip(n14793), .ck(clk), .q(\LUT[82][15] ) );
  dp_1 \LUT_reg[82][14]  ( .ip(n14792), .ck(clk), .q(\LUT[82][14] ) );
  dp_1 \LUT_reg[82][13]  ( .ip(n14791), .ck(clk), .q(\LUT[82][13] ) );
  dp_1 \LUT_reg[82][12]  ( .ip(n14790), .ck(clk), .q(\LUT[82][12] ) );
  dp_1 \LUT_reg[82][11]  ( .ip(n14789), .ck(clk), .q(\LUT[82][11] ) );
  dp_1 \LUT_reg[82][10]  ( .ip(n14788), .ck(clk), .q(\LUT[82][10] ) );
  dp_1 \LUT_reg[82][9]  ( .ip(n14787), .ck(clk), .q(\LUT[82][9] ) );
  dp_1 \LUT_reg[82][8]  ( .ip(n14786), .ck(clk), .q(\LUT[82][8] ) );
  dp_1 \LUT_reg[82][7]  ( .ip(n14785), .ck(clk), .q(\LUT[82][7] ) );
  dp_1 \LUT_reg[82][6]  ( .ip(n14784), .ck(clk), .q(\LUT[82][6] ) );
  dp_1 \LUT_reg[82][5]  ( .ip(n14783), .ck(clk), .q(\LUT[82][5] ) );
  dp_1 \LUT_reg[82][4]  ( .ip(n14782), .ck(clk), .q(\LUT[82][4] ) );
  dp_1 \LUT_reg[82][3]  ( .ip(n14781), .ck(clk), .q(\LUT[82][3] ) );
  dp_1 \LUT_reg[82][2]  ( .ip(n14780), .ck(clk), .q(\LUT[82][2] ) );
  dp_1 \LUT_reg[82][1]  ( .ip(n14779), .ck(clk), .q(\LUT[82][1] ) );
  dp_1 \LUT_reg[82][0]  ( .ip(n14778), .ck(clk), .q(\LUT[82][0] ) );
  dp_1 \LUT_reg[81][15]  ( .ip(n14777), .ck(clk), .q(\LUT[81][15] ) );
  dp_1 \LUT_reg[81][14]  ( .ip(n14776), .ck(clk), .q(\LUT[81][14] ) );
  dp_1 \LUT_reg[81][13]  ( .ip(n14775), .ck(clk), .q(\LUT[81][13] ) );
  dp_1 \LUT_reg[81][12]  ( .ip(n14774), .ck(clk), .q(\LUT[81][12] ) );
  dp_1 \LUT_reg[81][11]  ( .ip(n14773), .ck(clk), .q(\LUT[81][11] ) );
  dp_1 \LUT_reg[81][10]  ( .ip(n14772), .ck(clk), .q(\LUT[81][10] ) );
  dp_1 \LUT_reg[81][9]  ( .ip(n14771), .ck(clk), .q(\LUT[81][9] ) );
  dp_1 \LUT_reg[81][8]  ( .ip(n14770), .ck(clk), .q(\LUT[81][8] ) );
  dp_1 \LUT_reg[81][7]  ( .ip(n14769), .ck(clk), .q(\LUT[81][7] ) );
  dp_1 \LUT_reg[81][6]  ( .ip(n14768), .ck(clk), .q(\LUT[81][6] ) );
  dp_1 \LUT_reg[81][5]  ( .ip(n14767), .ck(clk), .q(\LUT[81][5] ) );
  dp_1 \LUT_reg[81][4]  ( .ip(n14766), .ck(clk), .q(\LUT[81][4] ) );
  dp_1 \LUT_reg[81][3]  ( .ip(n14765), .ck(clk), .q(\LUT[81][3] ) );
  dp_1 \LUT_reg[81][2]  ( .ip(n14764), .ck(clk), .q(\LUT[81][2] ) );
  dp_1 \LUT_reg[81][1]  ( .ip(n14763), .ck(clk), .q(\LUT[81][1] ) );
  dp_1 \LUT_reg[81][0]  ( .ip(n14762), .ck(clk), .q(\LUT[81][0] ) );
  dp_1 \LUT_reg[80][15]  ( .ip(n14761), .ck(clk), .q(\LUT[80][15] ) );
  dp_1 \LUT_reg[80][14]  ( .ip(n14760), .ck(clk), .q(\LUT[80][14] ) );
  dp_1 \LUT_reg[80][13]  ( .ip(n14759), .ck(clk), .q(\LUT[80][13] ) );
  dp_1 \LUT_reg[80][12]  ( .ip(n14758), .ck(clk), .q(\LUT[80][12] ) );
  dp_1 \LUT_reg[80][11]  ( .ip(n14757), .ck(clk), .q(\LUT[80][11] ) );
  dp_1 \LUT_reg[80][10]  ( .ip(n14756), .ck(clk), .q(\LUT[80][10] ) );
  dp_1 \LUT_reg[80][9]  ( .ip(n14755), .ck(clk), .q(\LUT[80][9] ) );
  dp_1 \LUT_reg[80][8]  ( .ip(n14754), .ck(clk), .q(\LUT[80][8] ) );
  dp_1 \LUT_reg[80][7]  ( .ip(n14753), .ck(clk), .q(\LUT[80][7] ) );
  dp_1 \LUT_reg[80][6]  ( .ip(n14752), .ck(clk), .q(\LUT[80][6] ) );
  dp_1 \LUT_reg[80][5]  ( .ip(n14751), .ck(clk), .q(\LUT[80][5] ) );
  dp_1 \LUT_reg[80][4]  ( .ip(n14750), .ck(clk), .q(\LUT[80][4] ) );
  dp_1 \LUT_reg[80][3]  ( .ip(n14749), .ck(clk), .q(\LUT[80][3] ) );
  dp_1 \LUT_reg[80][2]  ( .ip(n14748), .ck(clk), .q(\LUT[80][2] ) );
  dp_1 \LUT_reg[80][1]  ( .ip(n14747), .ck(clk), .q(\LUT[80][1] ) );
  dp_1 \LUT_reg[80][0]  ( .ip(n14746), .ck(clk), .q(\LUT[80][0] ) );
  dp_1 \LUT_reg[79][15]  ( .ip(n14745), .ck(clk), .q(\LUT[79][15] ) );
  dp_1 \LUT_reg[79][14]  ( .ip(n14744), .ck(clk), .q(\LUT[79][14] ) );
  dp_1 \LUT_reg[79][13]  ( .ip(n14743), .ck(clk), .q(\LUT[79][13] ) );
  dp_1 \LUT_reg[79][12]  ( .ip(n14742), .ck(clk), .q(\LUT[79][12] ) );
  dp_1 \LUT_reg[79][11]  ( .ip(n14741), .ck(clk), .q(\LUT[79][11] ) );
  dp_1 \LUT_reg[79][10]  ( .ip(n14740), .ck(clk), .q(\LUT[79][10] ) );
  dp_1 \LUT_reg[79][9]  ( .ip(n14739), .ck(clk), .q(\LUT[79][9] ) );
  dp_1 \LUT_reg[79][8]  ( .ip(n14738), .ck(clk), .q(\LUT[79][8] ) );
  dp_1 \LUT_reg[79][7]  ( .ip(n14737), .ck(clk), .q(\LUT[79][7] ) );
  dp_1 \LUT_reg[79][6]  ( .ip(n14736), .ck(clk), .q(\LUT[79][6] ) );
  dp_1 \LUT_reg[79][5]  ( .ip(n14735), .ck(clk), .q(\LUT[79][5] ) );
  dp_1 \LUT_reg[79][4]  ( .ip(n14734), .ck(clk), .q(\LUT[79][4] ) );
  dp_1 \LUT_reg[79][3]  ( .ip(n14733), .ck(clk), .q(\LUT[79][3] ) );
  dp_1 \LUT_reg[79][2]  ( .ip(n14732), .ck(clk), .q(\LUT[79][2] ) );
  dp_1 \LUT_reg[79][1]  ( .ip(n14731), .ck(clk), .q(\LUT[79][1] ) );
  dp_1 \LUT_reg[79][0]  ( .ip(n14730), .ck(clk), .q(\LUT[79][0] ) );
  dp_1 \LUT_reg[78][15]  ( .ip(n14729), .ck(clk), .q(\LUT[78][15] ) );
  dp_1 \LUT_reg[78][14]  ( .ip(n14728), .ck(clk), .q(\LUT[78][14] ) );
  dp_1 \LUT_reg[78][13]  ( .ip(n14727), .ck(clk), .q(\LUT[78][13] ) );
  dp_1 \LUT_reg[78][12]  ( .ip(n14726), .ck(clk), .q(\LUT[78][12] ) );
  dp_1 \LUT_reg[78][11]  ( .ip(n14725), .ck(clk), .q(\LUT[78][11] ) );
  dp_1 \LUT_reg[78][10]  ( .ip(n14724), .ck(clk), .q(\LUT[78][10] ) );
  dp_1 \LUT_reg[78][9]  ( .ip(n14723), .ck(clk), .q(\LUT[78][9] ) );
  dp_1 \LUT_reg[78][8]  ( .ip(n14722), .ck(clk), .q(\LUT[78][8] ) );
  dp_1 \LUT_reg[78][7]  ( .ip(n14721), .ck(clk), .q(\LUT[78][7] ) );
  dp_1 \LUT_reg[78][6]  ( .ip(n14720), .ck(clk), .q(\LUT[78][6] ) );
  dp_1 \LUT_reg[78][5]  ( .ip(n14719), .ck(clk), .q(\LUT[78][5] ) );
  dp_1 \LUT_reg[78][4]  ( .ip(n14718), .ck(clk), .q(\LUT[78][4] ) );
  dp_1 \LUT_reg[78][3]  ( .ip(n14717), .ck(clk), .q(\LUT[78][3] ) );
  dp_1 \LUT_reg[78][2]  ( .ip(n14716), .ck(clk), .q(\LUT[78][2] ) );
  dp_1 \LUT_reg[78][1]  ( .ip(n14715), .ck(clk), .q(\LUT[78][1] ) );
  dp_1 \LUT_reg[78][0]  ( .ip(n14714), .ck(clk), .q(\LUT[78][0] ) );
  dp_1 \LUT_reg[77][15]  ( .ip(n14713), .ck(clk), .q(\LUT[77][15] ) );
  dp_1 \LUT_reg[77][14]  ( .ip(n14712), .ck(clk), .q(\LUT[77][14] ) );
  dp_1 \LUT_reg[77][13]  ( .ip(n14711), .ck(clk), .q(\LUT[77][13] ) );
  dp_1 \LUT_reg[77][12]  ( .ip(n14710), .ck(clk), .q(\LUT[77][12] ) );
  dp_1 \LUT_reg[77][11]  ( .ip(n14709), .ck(clk), .q(\LUT[77][11] ) );
  dp_1 \LUT_reg[77][10]  ( .ip(n14708), .ck(clk), .q(\LUT[77][10] ) );
  dp_1 \LUT_reg[77][9]  ( .ip(n14707), .ck(clk), .q(\LUT[77][9] ) );
  dp_1 \LUT_reg[77][8]  ( .ip(n14706), .ck(clk), .q(\LUT[77][8] ) );
  dp_1 \LUT_reg[77][7]  ( .ip(n14705), .ck(clk), .q(\LUT[77][7] ) );
  dp_1 \LUT_reg[77][6]  ( .ip(n14704), .ck(clk), .q(\LUT[77][6] ) );
  dp_1 \LUT_reg[77][5]  ( .ip(n14703), .ck(clk), .q(\LUT[77][5] ) );
  dp_1 \LUT_reg[77][4]  ( .ip(n14702), .ck(clk), .q(\LUT[77][4] ) );
  dp_1 \LUT_reg[77][3]  ( .ip(n14701), .ck(clk), .q(\LUT[77][3] ) );
  dp_1 \LUT_reg[77][2]  ( .ip(n14700), .ck(clk), .q(\LUT[77][2] ) );
  dp_1 \LUT_reg[77][1]  ( .ip(n14699), .ck(clk), .q(\LUT[77][1] ) );
  dp_1 \LUT_reg[77][0]  ( .ip(n14698), .ck(clk), .q(\LUT[77][0] ) );
  dp_1 \LUT_reg[76][15]  ( .ip(n14697), .ck(clk), .q(\LUT[76][15] ) );
  dp_1 \LUT_reg[76][14]  ( .ip(n14696), .ck(clk), .q(\LUT[76][14] ) );
  dp_1 \LUT_reg[76][13]  ( .ip(n14695), .ck(clk), .q(\LUT[76][13] ) );
  dp_1 \LUT_reg[76][12]  ( .ip(n14694), .ck(clk), .q(\LUT[76][12] ) );
  dp_1 \LUT_reg[76][11]  ( .ip(n14693), .ck(clk), .q(\LUT[76][11] ) );
  dp_1 \LUT_reg[76][10]  ( .ip(n14692), .ck(clk), .q(\LUT[76][10] ) );
  dp_1 \LUT_reg[76][9]  ( .ip(n14691), .ck(clk), .q(\LUT[76][9] ) );
  dp_1 \LUT_reg[76][8]  ( .ip(n14690), .ck(clk), .q(\LUT[76][8] ) );
  dp_1 \LUT_reg[76][7]  ( .ip(n14689), .ck(clk), .q(\LUT[76][7] ) );
  dp_1 \LUT_reg[76][6]  ( .ip(n14688), .ck(clk), .q(\LUT[76][6] ) );
  dp_1 \LUT_reg[76][5]  ( .ip(n14687), .ck(clk), .q(\LUT[76][5] ) );
  dp_1 \LUT_reg[76][4]  ( .ip(n14686), .ck(clk), .q(\LUT[76][4] ) );
  dp_1 \LUT_reg[76][3]  ( .ip(n14685), .ck(clk), .q(\LUT[76][3] ) );
  dp_1 \LUT_reg[76][2]  ( .ip(n14684), .ck(clk), .q(\LUT[76][2] ) );
  dp_1 \LUT_reg[76][1]  ( .ip(n14683), .ck(clk), .q(\LUT[76][1] ) );
  dp_1 \LUT_reg[76][0]  ( .ip(n14682), .ck(clk), .q(\LUT[76][0] ) );
  dp_1 \LUT_reg[75][15]  ( .ip(n14681), .ck(clk), .q(\LUT[75][15] ) );
  dp_1 \LUT_reg[75][14]  ( .ip(n14680), .ck(clk), .q(\LUT[75][14] ) );
  dp_1 \LUT_reg[75][13]  ( .ip(n14679), .ck(clk), .q(\LUT[75][13] ) );
  dp_1 \LUT_reg[75][12]  ( .ip(n14678), .ck(clk), .q(\LUT[75][12] ) );
  dp_1 \LUT_reg[75][11]  ( .ip(n14677), .ck(clk), .q(\LUT[75][11] ) );
  dp_1 \LUT_reg[75][10]  ( .ip(n14676), .ck(clk), .q(\LUT[75][10] ) );
  dp_1 \LUT_reg[75][9]  ( .ip(n14675), .ck(clk), .q(\LUT[75][9] ) );
  dp_1 \LUT_reg[75][8]  ( .ip(n14674), .ck(clk), .q(\LUT[75][8] ) );
  dp_1 \LUT_reg[75][7]  ( .ip(n14673), .ck(clk), .q(\LUT[75][7] ) );
  dp_1 \LUT_reg[75][6]  ( .ip(n14672), .ck(clk), .q(\LUT[75][6] ) );
  dp_1 \LUT_reg[75][5]  ( .ip(n14671), .ck(clk), .q(\LUT[75][5] ) );
  dp_1 \LUT_reg[75][4]  ( .ip(n14670), .ck(clk), .q(\LUT[75][4] ) );
  dp_1 \LUT_reg[75][3]  ( .ip(n14669), .ck(clk), .q(\LUT[75][3] ) );
  dp_1 \LUT_reg[75][2]  ( .ip(n14668), .ck(clk), .q(\LUT[75][2] ) );
  dp_1 \LUT_reg[75][1]  ( .ip(n14667), .ck(clk), .q(\LUT[75][1] ) );
  dp_1 \LUT_reg[75][0]  ( .ip(n14666), .ck(clk), .q(\LUT[75][0] ) );
  dp_1 \LUT_reg[74][15]  ( .ip(n14665), .ck(clk), .q(\LUT[74][15] ) );
  dp_1 \LUT_reg[74][14]  ( .ip(n14664), .ck(clk), .q(\LUT[74][14] ) );
  dp_1 \LUT_reg[74][13]  ( .ip(n14663), .ck(clk), .q(\LUT[74][13] ) );
  dp_1 \LUT_reg[74][12]  ( .ip(n14662), .ck(clk), .q(\LUT[74][12] ) );
  dp_1 \LUT_reg[74][11]  ( .ip(n14661), .ck(clk), .q(\LUT[74][11] ) );
  dp_1 \LUT_reg[74][10]  ( .ip(n14660), .ck(clk), .q(\LUT[74][10] ) );
  dp_1 \LUT_reg[74][9]  ( .ip(n14659), .ck(clk), .q(\LUT[74][9] ) );
  dp_1 \LUT_reg[74][8]  ( .ip(n14658), .ck(clk), .q(\LUT[74][8] ) );
  dp_1 \LUT_reg[74][7]  ( .ip(n14657), .ck(clk), .q(\LUT[74][7] ) );
  dp_1 \LUT_reg[74][6]  ( .ip(n14656), .ck(clk), .q(\LUT[74][6] ) );
  dp_1 \LUT_reg[74][5]  ( .ip(n14655), .ck(clk), .q(\LUT[74][5] ) );
  dp_1 \LUT_reg[74][4]  ( .ip(n14654), .ck(clk), .q(\LUT[74][4] ) );
  dp_1 \LUT_reg[74][3]  ( .ip(n14653), .ck(clk), .q(\LUT[74][3] ) );
  dp_1 \LUT_reg[74][2]  ( .ip(n14652), .ck(clk), .q(\LUT[74][2] ) );
  dp_1 \LUT_reg[74][1]  ( .ip(n14651), .ck(clk), .q(\LUT[74][1] ) );
  dp_1 \LUT_reg[74][0]  ( .ip(n14650), .ck(clk), .q(\LUT[74][0] ) );
  dp_1 \LUT_reg[73][15]  ( .ip(n14649), .ck(clk), .q(\LUT[73][15] ) );
  dp_1 \LUT_reg[73][14]  ( .ip(n14648), .ck(clk), .q(\LUT[73][14] ) );
  dp_1 \LUT_reg[73][13]  ( .ip(n14647), .ck(clk), .q(\LUT[73][13] ) );
  dp_1 \LUT_reg[73][12]  ( .ip(n14646), .ck(clk), .q(\LUT[73][12] ) );
  dp_1 \LUT_reg[73][11]  ( .ip(n14645), .ck(clk), .q(\LUT[73][11] ) );
  dp_1 \LUT_reg[73][10]  ( .ip(n14644), .ck(clk), .q(\LUT[73][10] ) );
  dp_1 \LUT_reg[73][9]  ( .ip(n14643), .ck(clk), .q(\LUT[73][9] ) );
  dp_1 \LUT_reg[73][8]  ( .ip(n14642), .ck(clk), .q(\LUT[73][8] ) );
  dp_1 \LUT_reg[73][7]  ( .ip(n14641), .ck(clk), .q(\LUT[73][7] ) );
  dp_1 \LUT_reg[73][6]  ( .ip(n14640), .ck(clk), .q(\LUT[73][6] ) );
  dp_1 \LUT_reg[73][5]  ( .ip(n14639), .ck(clk), .q(\LUT[73][5] ) );
  dp_1 \LUT_reg[73][4]  ( .ip(n14638), .ck(clk), .q(\LUT[73][4] ) );
  dp_1 \LUT_reg[73][3]  ( .ip(n14637), .ck(clk), .q(\LUT[73][3] ) );
  dp_1 \LUT_reg[73][2]  ( .ip(n14636), .ck(clk), .q(\LUT[73][2] ) );
  dp_1 \LUT_reg[73][1]  ( .ip(n14635), .ck(clk), .q(\LUT[73][1] ) );
  dp_1 \LUT_reg[73][0]  ( .ip(n14634), .ck(clk), .q(\LUT[73][0] ) );
  dp_1 \LUT_reg[72][15]  ( .ip(n14633), .ck(clk), .q(\LUT[72][15] ) );
  dp_1 \LUT_reg[72][14]  ( .ip(n14632), .ck(clk), .q(\LUT[72][14] ) );
  dp_1 \LUT_reg[72][13]  ( .ip(n14631), .ck(clk), .q(\LUT[72][13] ) );
  dp_1 \LUT_reg[72][12]  ( .ip(n14630), .ck(clk), .q(\LUT[72][12] ) );
  dp_1 \LUT_reg[72][11]  ( .ip(n14629), .ck(clk), .q(\LUT[72][11] ) );
  dp_1 \LUT_reg[72][10]  ( .ip(n14628), .ck(clk), .q(\LUT[72][10] ) );
  dp_1 \LUT_reg[72][9]  ( .ip(n14627), .ck(clk), .q(\LUT[72][9] ) );
  dp_1 \LUT_reg[72][8]  ( .ip(n14626), .ck(clk), .q(\LUT[72][8] ) );
  dp_1 \LUT_reg[72][7]  ( .ip(n14625), .ck(clk), .q(\LUT[72][7] ) );
  dp_1 \LUT_reg[72][6]  ( .ip(n14624), .ck(clk), .q(\LUT[72][6] ) );
  dp_1 \LUT_reg[72][5]  ( .ip(n14623), .ck(clk), .q(\LUT[72][5] ) );
  dp_1 \LUT_reg[72][4]  ( .ip(n14622), .ck(clk), .q(\LUT[72][4] ) );
  dp_1 \LUT_reg[72][3]  ( .ip(n14621), .ck(clk), .q(\LUT[72][3] ) );
  dp_1 \LUT_reg[72][2]  ( .ip(n14620), .ck(clk), .q(\LUT[72][2] ) );
  dp_1 \LUT_reg[72][1]  ( .ip(n14619), .ck(clk), .q(\LUT[72][1] ) );
  dp_1 \LUT_reg[72][0]  ( .ip(n14618), .ck(clk), .q(\LUT[72][0] ) );
  dp_1 \LUT_reg[71][15]  ( .ip(n14617), .ck(clk), .q(\LUT[71][15] ) );
  dp_1 \LUT_reg[71][14]  ( .ip(n14616), .ck(clk), .q(\LUT[71][14] ) );
  dp_1 \LUT_reg[71][13]  ( .ip(n14615), .ck(clk), .q(\LUT[71][13] ) );
  dp_1 \LUT_reg[71][12]  ( .ip(n14614), .ck(clk), .q(\LUT[71][12] ) );
  dp_1 \LUT_reg[71][11]  ( .ip(n14613), .ck(clk), .q(\LUT[71][11] ) );
  dp_1 \LUT_reg[71][10]  ( .ip(n14612), .ck(clk), .q(\LUT[71][10] ) );
  dp_1 \LUT_reg[71][9]  ( .ip(n14611), .ck(clk), .q(\LUT[71][9] ) );
  dp_1 \LUT_reg[71][8]  ( .ip(n14610), .ck(clk), .q(\LUT[71][8] ) );
  dp_1 \LUT_reg[71][7]  ( .ip(n14609), .ck(clk), .q(\LUT[71][7] ) );
  dp_1 \LUT_reg[71][6]  ( .ip(n14608), .ck(clk), .q(\LUT[71][6] ) );
  dp_1 \LUT_reg[71][5]  ( .ip(n14607), .ck(clk), .q(\LUT[71][5] ) );
  dp_1 \LUT_reg[71][4]  ( .ip(n14606), .ck(clk), .q(\LUT[71][4] ) );
  dp_1 \LUT_reg[71][3]  ( .ip(n14605), .ck(clk), .q(\LUT[71][3] ) );
  dp_1 \LUT_reg[71][2]  ( .ip(n14604), .ck(clk), .q(\LUT[71][2] ) );
  dp_1 \LUT_reg[71][1]  ( .ip(n14603), .ck(clk), .q(\LUT[71][1] ) );
  dp_1 \LUT_reg[71][0]  ( .ip(n14602), .ck(clk), .q(\LUT[71][0] ) );
  dp_1 \LUT_reg[70][15]  ( .ip(n14601), .ck(clk), .q(\LUT[70][15] ) );
  dp_1 \LUT_reg[70][14]  ( .ip(n14600), .ck(clk), .q(\LUT[70][14] ) );
  dp_1 \LUT_reg[70][13]  ( .ip(n14599), .ck(clk), .q(\LUT[70][13] ) );
  dp_1 \LUT_reg[70][12]  ( .ip(n14598), .ck(clk), .q(\LUT[70][12] ) );
  dp_1 \LUT_reg[70][11]  ( .ip(n14597), .ck(clk), .q(\LUT[70][11] ) );
  dp_1 \LUT_reg[70][10]  ( .ip(n14596), .ck(clk), .q(\LUT[70][10] ) );
  dp_1 \LUT_reg[70][9]  ( .ip(n14595), .ck(clk), .q(\LUT[70][9] ) );
  dp_1 \LUT_reg[70][8]  ( .ip(n14594), .ck(clk), .q(\LUT[70][8] ) );
  dp_1 \LUT_reg[70][7]  ( .ip(n14593), .ck(clk), .q(\LUT[70][7] ) );
  dp_1 \LUT_reg[70][6]  ( .ip(n14592), .ck(clk), .q(\LUT[70][6] ) );
  dp_1 \LUT_reg[70][5]  ( .ip(n14591), .ck(clk), .q(\LUT[70][5] ) );
  dp_1 \LUT_reg[70][4]  ( .ip(n14590), .ck(clk), .q(\LUT[70][4] ) );
  dp_1 \LUT_reg[70][3]  ( .ip(n14589), .ck(clk), .q(\LUT[70][3] ) );
  dp_1 \LUT_reg[70][2]  ( .ip(n14588), .ck(clk), .q(\LUT[70][2] ) );
  dp_1 \LUT_reg[70][1]  ( .ip(n14587), .ck(clk), .q(\LUT[70][1] ) );
  dp_1 \LUT_reg[70][0]  ( .ip(n14586), .ck(clk), .q(\LUT[70][0] ) );
  dp_1 \LUT_reg[69][15]  ( .ip(n14585), .ck(clk), .q(\LUT[69][15] ) );
  dp_1 \LUT_reg[69][14]  ( .ip(n14584), .ck(clk), .q(\LUT[69][14] ) );
  dp_1 \LUT_reg[69][13]  ( .ip(n14583), .ck(clk), .q(\LUT[69][13] ) );
  dp_1 \LUT_reg[69][12]  ( .ip(n14582), .ck(clk), .q(\LUT[69][12] ) );
  dp_1 \LUT_reg[69][11]  ( .ip(n14581), .ck(clk), .q(\LUT[69][11] ) );
  dp_1 \LUT_reg[69][10]  ( .ip(n14580), .ck(clk), .q(\LUT[69][10] ) );
  dp_1 \LUT_reg[69][9]  ( .ip(n14579), .ck(clk), .q(\LUT[69][9] ) );
  dp_1 \LUT_reg[69][8]  ( .ip(n14578), .ck(clk), .q(\LUT[69][8] ) );
  dp_1 \LUT_reg[69][7]  ( .ip(n14577), .ck(clk), .q(\LUT[69][7] ) );
  dp_1 \LUT_reg[69][6]  ( .ip(n14576), .ck(clk), .q(\LUT[69][6] ) );
  dp_1 \LUT_reg[69][5]  ( .ip(n14575), .ck(clk), .q(\LUT[69][5] ) );
  dp_1 \LUT_reg[69][4]  ( .ip(n14574), .ck(clk), .q(\LUT[69][4] ) );
  dp_1 \LUT_reg[69][3]  ( .ip(n14573), .ck(clk), .q(\LUT[69][3] ) );
  dp_1 \LUT_reg[69][2]  ( .ip(n14572), .ck(clk), .q(\LUT[69][2] ) );
  dp_1 \LUT_reg[69][1]  ( .ip(n14571), .ck(clk), .q(\LUT[69][1] ) );
  dp_1 \LUT_reg[69][0]  ( .ip(n14570), .ck(clk), .q(\LUT[69][0] ) );
  dp_1 \LUT_reg[68][15]  ( .ip(n14569), .ck(clk), .q(\LUT[68][15] ) );
  dp_1 \LUT_reg[68][14]  ( .ip(n14568), .ck(clk), .q(\LUT[68][14] ) );
  dp_1 \LUT_reg[68][13]  ( .ip(n14567), .ck(clk), .q(\LUT[68][13] ) );
  dp_1 \LUT_reg[68][12]  ( .ip(n14566), .ck(clk), .q(\LUT[68][12] ) );
  dp_1 \LUT_reg[68][11]  ( .ip(n14565), .ck(clk), .q(\LUT[68][11] ) );
  dp_1 \LUT_reg[68][10]  ( .ip(n14564), .ck(clk), .q(\LUT[68][10] ) );
  dp_1 \LUT_reg[68][9]  ( .ip(n14563), .ck(clk), .q(\LUT[68][9] ) );
  dp_1 \LUT_reg[68][8]  ( .ip(n14562), .ck(clk), .q(\LUT[68][8] ) );
  dp_1 \LUT_reg[68][7]  ( .ip(n14561), .ck(clk), .q(\LUT[68][7] ) );
  dp_1 \LUT_reg[68][6]  ( .ip(n14560), .ck(clk), .q(\LUT[68][6] ) );
  dp_1 \LUT_reg[68][5]  ( .ip(n14559), .ck(clk), .q(\LUT[68][5] ) );
  dp_1 \LUT_reg[68][4]  ( .ip(n14558), .ck(clk), .q(\LUT[68][4] ) );
  dp_1 \LUT_reg[68][3]  ( .ip(n14557), .ck(clk), .q(\LUT[68][3] ) );
  dp_1 \LUT_reg[68][2]  ( .ip(n14556), .ck(clk), .q(\LUT[68][2] ) );
  dp_1 \LUT_reg[68][1]  ( .ip(n14555), .ck(clk), .q(\LUT[68][1] ) );
  dp_1 \LUT_reg[68][0]  ( .ip(n14554), .ck(clk), .q(\LUT[68][0] ) );
  dp_1 \LUT_reg[67][15]  ( .ip(n14553), .ck(clk), .q(\LUT[67][15] ) );
  dp_1 \LUT_reg[67][14]  ( .ip(n14552), .ck(clk), .q(\LUT[67][14] ) );
  dp_1 \LUT_reg[67][13]  ( .ip(n14551), .ck(clk), .q(\LUT[67][13] ) );
  dp_1 \LUT_reg[67][12]  ( .ip(n14550), .ck(clk), .q(\LUT[67][12] ) );
  dp_1 \LUT_reg[67][11]  ( .ip(n14549), .ck(clk), .q(\LUT[67][11] ) );
  dp_1 \LUT_reg[67][10]  ( .ip(n14548), .ck(clk), .q(\LUT[67][10] ) );
  dp_1 \LUT_reg[67][9]  ( .ip(n14547), .ck(clk), .q(\LUT[67][9] ) );
  dp_1 \LUT_reg[67][8]  ( .ip(n14546), .ck(clk), .q(\LUT[67][8] ) );
  dp_1 \LUT_reg[67][7]  ( .ip(n14545), .ck(clk), .q(\LUT[67][7] ) );
  dp_1 \LUT_reg[67][6]  ( .ip(n14544), .ck(clk), .q(\LUT[67][6] ) );
  dp_1 \LUT_reg[67][5]  ( .ip(n14543), .ck(clk), .q(\LUT[67][5] ) );
  dp_1 \LUT_reg[67][4]  ( .ip(n14542), .ck(clk), .q(\LUT[67][4] ) );
  dp_1 \LUT_reg[67][3]  ( .ip(n14541), .ck(clk), .q(\LUT[67][3] ) );
  dp_1 \LUT_reg[67][2]  ( .ip(n14540), .ck(clk), .q(\LUT[67][2] ) );
  dp_1 \LUT_reg[67][1]  ( .ip(n14539), .ck(clk), .q(\LUT[67][1] ) );
  dp_1 \LUT_reg[67][0]  ( .ip(n14538), .ck(clk), .q(\LUT[67][0] ) );
  dp_1 \LUT_reg[66][15]  ( .ip(n14537), .ck(clk), .q(\LUT[66][15] ) );
  dp_1 \LUT_reg[66][14]  ( .ip(n14536), .ck(clk), .q(\LUT[66][14] ) );
  dp_1 \LUT_reg[66][13]  ( .ip(n14535), .ck(clk), .q(\LUT[66][13] ) );
  dp_1 \LUT_reg[66][12]  ( .ip(n14534), .ck(clk), .q(\LUT[66][12] ) );
  dp_1 \LUT_reg[66][11]  ( .ip(n14533), .ck(clk), .q(\LUT[66][11] ) );
  dp_1 \LUT_reg[66][10]  ( .ip(n14532), .ck(clk), .q(\LUT[66][10] ) );
  dp_1 \LUT_reg[66][9]  ( .ip(n14531), .ck(clk), .q(\LUT[66][9] ) );
  dp_1 \LUT_reg[66][8]  ( .ip(n14530), .ck(clk), .q(\LUT[66][8] ) );
  dp_1 \LUT_reg[66][7]  ( .ip(n14529), .ck(clk), .q(\LUT[66][7] ) );
  dp_1 \LUT_reg[66][6]  ( .ip(n14528), .ck(clk), .q(\LUT[66][6] ) );
  dp_1 \LUT_reg[66][5]  ( .ip(n14527), .ck(clk), .q(\LUT[66][5] ) );
  dp_1 \LUT_reg[66][4]  ( .ip(n14526), .ck(clk), .q(\LUT[66][4] ) );
  dp_1 \LUT_reg[66][3]  ( .ip(n14525), .ck(clk), .q(\LUT[66][3] ) );
  dp_1 \LUT_reg[66][2]  ( .ip(n14524), .ck(clk), .q(\LUT[66][2] ) );
  dp_1 \LUT_reg[66][1]  ( .ip(n14523), .ck(clk), .q(\LUT[66][1] ) );
  dp_1 \LUT_reg[66][0]  ( .ip(n14522), .ck(clk), .q(\LUT[66][0] ) );
  dp_1 \LUT_reg[65][15]  ( .ip(n14521), .ck(clk), .q(\LUT[65][15] ) );
  dp_1 \LUT_reg[65][14]  ( .ip(n14520), .ck(clk), .q(\LUT[65][14] ) );
  dp_1 \LUT_reg[65][13]  ( .ip(n14519), .ck(clk), .q(\LUT[65][13] ) );
  dp_1 \LUT_reg[65][12]  ( .ip(n14518), .ck(clk), .q(\LUT[65][12] ) );
  dp_1 \LUT_reg[65][11]  ( .ip(n14517), .ck(clk), .q(\LUT[65][11] ) );
  dp_1 \LUT_reg[65][10]  ( .ip(n14516), .ck(clk), .q(\LUT[65][10] ) );
  dp_1 \LUT_reg[65][9]  ( .ip(n14515), .ck(clk), .q(\LUT[65][9] ) );
  dp_1 \LUT_reg[65][8]  ( .ip(n14514), .ck(clk), .q(\LUT[65][8] ) );
  dp_1 \LUT_reg[65][7]  ( .ip(n14513), .ck(clk), .q(\LUT[65][7] ) );
  dp_1 \LUT_reg[65][6]  ( .ip(n14512), .ck(clk), .q(\LUT[65][6] ) );
  dp_1 \LUT_reg[65][5]  ( .ip(n14511), .ck(clk), .q(\LUT[65][5] ) );
  dp_1 \LUT_reg[65][4]  ( .ip(n14510), .ck(clk), .q(\LUT[65][4] ) );
  dp_1 \LUT_reg[65][3]  ( .ip(n14509), .ck(clk), .q(\LUT[65][3] ) );
  dp_1 \LUT_reg[65][2]  ( .ip(n14508), .ck(clk), .q(\LUT[65][2] ) );
  dp_1 \LUT_reg[65][1]  ( .ip(n14507), .ck(clk), .q(\LUT[65][1] ) );
  dp_1 \LUT_reg[65][0]  ( .ip(n14506), .ck(clk), .q(\LUT[65][0] ) );
  dp_1 \LUT_reg[64][15]  ( .ip(n14505), .ck(clk), .q(\LUT[64][15] ) );
  dp_1 \LUT_reg[64][14]  ( .ip(n14504), .ck(clk), .q(\LUT[64][14] ) );
  dp_1 \LUT_reg[64][13]  ( .ip(n14503), .ck(clk), .q(\LUT[64][13] ) );
  dp_1 \LUT_reg[64][12]  ( .ip(n14502), .ck(clk), .q(\LUT[64][12] ) );
  dp_1 \LUT_reg[64][11]  ( .ip(n14501), .ck(clk), .q(\LUT[64][11] ) );
  dp_1 \LUT_reg[64][10]  ( .ip(n14500), .ck(clk), .q(\LUT[64][10] ) );
  dp_1 \LUT_reg[64][9]  ( .ip(n14499), .ck(clk), .q(\LUT[64][9] ) );
  dp_1 \LUT_reg[64][8]  ( .ip(n14498), .ck(clk), .q(\LUT[64][8] ) );
  dp_1 \LUT_reg[64][7]  ( .ip(n14497), .ck(clk), .q(\LUT[64][7] ) );
  dp_1 \LUT_reg[64][6]  ( .ip(n14496), .ck(clk), .q(\LUT[64][6] ) );
  dp_1 \LUT_reg[64][5]  ( .ip(n14495), .ck(clk), .q(\LUT[64][5] ) );
  dp_1 \LUT_reg[64][4]  ( .ip(n14494), .ck(clk), .q(\LUT[64][4] ) );
  dp_1 \LUT_reg[64][3]  ( .ip(n14493), .ck(clk), .q(\LUT[64][3] ) );
  dp_1 \LUT_reg[64][2]  ( .ip(n14492), .ck(clk), .q(\LUT[64][2] ) );
  dp_1 \LUT_reg[64][1]  ( .ip(n14491), .ck(clk), .q(\LUT[64][1] ) );
  dp_1 \LUT_reg[64][0]  ( .ip(n14490), .ck(clk), .q(\LUT[64][0] ) );
  dp_1 \LUT_reg[63][15]  ( .ip(n14489), .ck(clk), .q(\LUT[63][15] ) );
  dp_1 \LUT_reg[63][14]  ( .ip(n14488), .ck(clk), .q(\LUT[63][14] ) );
  dp_1 \LUT_reg[63][13]  ( .ip(n14487), .ck(clk), .q(\LUT[63][13] ) );
  dp_1 \LUT_reg[63][12]  ( .ip(n14486), .ck(clk), .q(\LUT[63][12] ) );
  dp_1 \LUT_reg[63][11]  ( .ip(n14485), .ck(clk), .q(\LUT[63][11] ) );
  dp_1 \LUT_reg[63][10]  ( .ip(n14484), .ck(clk), .q(\LUT[63][10] ) );
  dp_1 \LUT_reg[63][9]  ( .ip(n14483), .ck(clk), .q(\LUT[63][9] ) );
  dp_1 \LUT_reg[63][8]  ( .ip(n14482), .ck(clk), .q(\LUT[63][8] ) );
  dp_1 \LUT_reg[63][7]  ( .ip(n14481), .ck(clk), .q(\LUT[63][7] ) );
  dp_1 \LUT_reg[63][6]  ( .ip(n14480), .ck(clk), .q(\LUT[63][6] ) );
  dp_1 \LUT_reg[63][5]  ( .ip(n14479), .ck(clk), .q(\LUT[63][5] ) );
  dp_1 \LUT_reg[63][4]  ( .ip(n14478), .ck(clk), .q(\LUT[63][4] ) );
  dp_1 \LUT_reg[63][3]  ( .ip(n14477), .ck(clk), .q(\LUT[63][3] ) );
  dp_1 \LUT_reg[63][2]  ( .ip(n14476), .ck(clk), .q(\LUT[63][2] ) );
  dp_1 \LUT_reg[63][1]  ( .ip(n14475), .ck(clk), .q(\LUT[63][1] ) );
  dp_1 \LUT_reg[63][0]  ( .ip(n14474), .ck(clk), .q(\LUT[63][0] ) );
  dp_1 \LUT_reg[62][15]  ( .ip(n14473), .ck(clk), .q(\LUT[62][15] ) );
  dp_1 \LUT_reg[62][14]  ( .ip(n14472), .ck(clk), .q(\LUT[62][14] ) );
  dp_1 \LUT_reg[62][13]  ( .ip(n14471), .ck(clk), .q(\LUT[62][13] ) );
  dp_1 \LUT_reg[62][12]  ( .ip(n14470), .ck(clk), .q(\LUT[62][12] ) );
  dp_1 \LUT_reg[62][11]  ( .ip(n14469), .ck(clk), .q(\LUT[62][11] ) );
  dp_1 \LUT_reg[62][10]  ( .ip(n14468), .ck(clk), .q(\LUT[62][10] ) );
  dp_1 \LUT_reg[62][9]  ( .ip(n14467), .ck(clk), .q(\LUT[62][9] ) );
  dp_1 \LUT_reg[62][8]  ( .ip(n14466), .ck(clk), .q(\LUT[62][8] ) );
  dp_1 \LUT_reg[62][7]  ( .ip(n14465), .ck(clk), .q(\LUT[62][7] ) );
  dp_1 \LUT_reg[62][6]  ( .ip(n14464), .ck(clk), .q(\LUT[62][6] ) );
  dp_1 \LUT_reg[62][5]  ( .ip(n14463), .ck(clk), .q(\LUT[62][5] ) );
  dp_1 \LUT_reg[62][4]  ( .ip(n14462), .ck(clk), .q(\LUT[62][4] ) );
  dp_1 \LUT_reg[62][3]  ( .ip(n14461), .ck(clk), .q(\LUT[62][3] ) );
  dp_1 \LUT_reg[62][2]  ( .ip(n14460), .ck(clk), .q(\LUT[62][2] ) );
  dp_1 \LUT_reg[62][1]  ( .ip(n14459), .ck(clk), .q(\LUT[62][1] ) );
  dp_1 \LUT_reg[62][0]  ( .ip(n14458), .ck(clk), .q(\LUT[62][0] ) );
  dp_1 \LUT_reg[61][15]  ( .ip(n14457), .ck(clk), .q(\LUT[61][15] ) );
  dp_1 \LUT_reg[61][14]  ( .ip(n14456), .ck(clk), .q(\LUT[61][14] ) );
  dp_1 \LUT_reg[61][13]  ( .ip(n14455), .ck(clk), .q(\LUT[61][13] ) );
  dp_1 \LUT_reg[61][12]  ( .ip(n14454), .ck(clk), .q(\LUT[61][12] ) );
  dp_1 \LUT_reg[61][11]  ( .ip(n14453), .ck(clk), .q(\LUT[61][11] ) );
  dp_1 \LUT_reg[61][10]  ( .ip(n14452), .ck(clk), .q(\LUT[61][10] ) );
  dp_1 \LUT_reg[61][9]  ( .ip(n14451), .ck(clk), .q(\LUT[61][9] ) );
  dp_1 \LUT_reg[61][8]  ( .ip(n14450), .ck(clk), .q(\LUT[61][8] ) );
  dp_1 \LUT_reg[61][7]  ( .ip(n14449), .ck(clk), .q(\LUT[61][7] ) );
  dp_1 \LUT_reg[61][6]  ( .ip(n14448), .ck(clk), .q(\LUT[61][6] ) );
  dp_1 \LUT_reg[61][5]  ( .ip(n14447), .ck(clk), .q(\LUT[61][5] ) );
  dp_1 \LUT_reg[61][4]  ( .ip(n14446), .ck(clk), .q(\LUT[61][4] ) );
  dp_1 \LUT_reg[61][3]  ( .ip(n14445), .ck(clk), .q(\LUT[61][3] ) );
  dp_1 \LUT_reg[61][2]  ( .ip(n14444), .ck(clk), .q(\LUT[61][2] ) );
  dp_1 \LUT_reg[61][1]  ( .ip(n14443), .ck(clk), .q(\LUT[61][1] ) );
  dp_1 \LUT_reg[61][0]  ( .ip(n14442), .ck(clk), .q(\LUT[61][0] ) );
  dp_1 \LUT_reg[60][15]  ( .ip(n14441), .ck(clk), .q(\LUT[60][15] ) );
  dp_1 \LUT_reg[60][14]  ( .ip(n14440), .ck(clk), .q(\LUT[60][14] ) );
  dp_1 \LUT_reg[60][13]  ( .ip(n14439), .ck(clk), .q(\LUT[60][13] ) );
  dp_1 \LUT_reg[60][12]  ( .ip(n14438), .ck(clk), .q(\LUT[60][12] ) );
  dp_1 \LUT_reg[60][11]  ( .ip(n14437), .ck(clk), .q(\LUT[60][11] ) );
  dp_1 \LUT_reg[60][10]  ( .ip(n14436), .ck(clk), .q(\LUT[60][10] ) );
  dp_1 \LUT_reg[60][9]  ( .ip(n14435), .ck(clk), .q(\LUT[60][9] ) );
  dp_1 \LUT_reg[60][8]  ( .ip(n14434), .ck(clk), .q(\LUT[60][8] ) );
  dp_1 \LUT_reg[60][7]  ( .ip(n14433), .ck(clk), .q(\LUT[60][7] ) );
  dp_1 \LUT_reg[60][6]  ( .ip(n14432), .ck(clk), .q(\LUT[60][6] ) );
  dp_1 \LUT_reg[60][5]  ( .ip(n14431), .ck(clk), .q(\LUT[60][5] ) );
  dp_1 \LUT_reg[60][4]  ( .ip(n14430), .ck(clk), .q(\LUT[60][4] ) );
  dp_1 \LUT_reg[60][3]  ( .ip(n14429), .ck(clk), .q(\LUT[60][3] ) );
  dp_1 \LUT_reg[60][2]  ( .ip(n14428), .ck(clk), .q(\LUT[60][2] ) );
  dp_1 \LUT_reg[60][1]  ( .ip(n14427), .ck(clk), .q(\LUT[60][1] ) );
  dp_1 \LUT_reg[60][0]  ( .ip(n14426), .ck(clk), .q(\LUT[60][0] ) );
  dp_1 \LUT_reg[59][15]  ( .ip(n14425), .ck(clk), .q(\LUT[59][15] ) );
  dp_1 \LUT_reg[59][14]  ( .ip(n14424), .ck(clk), .q(\LUT[59][14] ) );
  dp_1 \LUT_reg[59][13]  ( .ip(n14423), .ck(clk), .q(\LUT[59][13] ) );
  dp_1 \LUT_reg[59][12]  ( .ip(n14422), .ck(clk), .q(\LUT[59][12] ) );
  dp_1 \LUT_reg[59][11]  ( .ip(n14421), .ck(clk), .q(\LUT[59][11] ) );
  dp_1 \LUT_reg[59][10]  ( .ip(n14420), .ck(clk), .q(\LUT[59][10] ) );
  dp_1 \LUT_reg[59][9]  ( .ip(n14419), .ck(clk), .q(\LUT[59][9] ) );
  dp_1 \LUT_reg[59][8]  ( .ip(n14418), .ck(clk), .q(\LUT[59][8] ) );
  dp_1 \LUT_reg[59][7]  ( .ip(n14417), .ck(clk), .q(\LUT[59][7] ) );
  dp_1 \LUT_reg[59][6]  ( .ip(n14416), .ck(clk), .q(\LUT[59][6] ) );
  dp_1 \LUT_reg[59][5]  ( .ip(n14415), .ck(clk), .q(\LUT[59][5] ) );
  dp_1 \LUT_reg[59][4]  ( .ip(n14414), .ck(clk), .q(\LUT[59][4] ) );
  dp_1 \LUT_reg[59][3]  ( .ip(n14413), .ck(clk), .q(\LUT[59][3] ) );
  dp_1 \LUT_reg[59][2]  ( .ip(n14412), .ck(clk), .q(\LUT[59][2] ) );
  dp_1 \LUT_reg[59][1]  ( .ip(n14411), .ck(clk), .q(\LUT[59][1] ) );
  dp_1 \LUT_reg[59][0]  ( .ip(n14410), .ck(clk), .q(\LUT[59][0] ) );
  dp_1 \LUT_reg[58][15]  ( .ip(n14409), .ck(clk), .q(\LUT[58][15] ) );
  dp_1 \LUT_reg[58][14]  ( .ip(n14408), .ck(clk), .q(\LUT[58][14] ) );
  dp_1 \LUT_reg[58][13]  ( .ip(n14407), .ck(clk), .q(\LUT[58][13] ) );
  dp_1 \LUT_reg[58][12]  ( .ip(n14406), .ck(clk), .q(\LUT[58][12] ) );
  dp_1 \LUT_reg[58][11]  ( .ip(n14405), .ck(clk), .q(\LUT[58][11] ) );
  dp_1 \LUT_reg[58][10]  ( .ip(n14404), .ck(clk), .q(\LUT[58][10] ) );
  dp_1 \LUT_reg[58][9]  ( .ip(n14403), .ck(clk), .q(\LUT[58][9] ) );
  dp_1 \LUT_reg[58][8]  ( .ip(n14402), .ck(clk), .q(\LUT[58][8] ) );
  dp_1 \LUT_reg[58][7]  ( .ip(n14401), .ck(clk), .q(\LUT[58][7] ) );
  dp_1 \LUT_reg[58][6]  ( .ip(n14400), .ck(clk), .q(\LUT[58][6] ) );
  dp_1 \LUT_reg[58][5]  ( .ip(n14399), .ck(clk), .q(\LUT[58][5] ) );
  dp_1 \LUT_reg[58][4]  ( .ip(n14398), .ck(clk), .q(\LUT[58][4] ) );
  dp_1 \LUT_reg[58][3]  ( .ip(n14397), .ck(clk), .q(\LUT[58][3] ) );
  dp_1 \LUT_reg[58][2]  ( .ip(n14396), .ck(clk), .q(\LUT[58][2] ) );
  dp_1 \LUT_reg[58][1]  ( .ip(n14395), .ck(clk), .q(\LUT[58][1] ) );
  dp_1 \LUT_reg[58][0]  ( .ip(n14394), .ck(clk), .q(\LUT[58][0] ) );
  dp_1 \LUT_reg[57][15]  ( .ip(n14393), .ck(clk), .q(\LUT[57][15] ) );
  dp_1 \LUT_reg[57][14]  ( .ip(n14392), .ck(clk), .q(\LUT[57][14] ) );
  dp_1 \LUT_reg[57][13]  ( .ip(n14391), .ck(clk), .q(\LUT[57][13] ) );
  dp_1 \LUT_reg[57][12]  ( .ip(n14390), .ck(clk), .q(\LUT[57][12] ) );
  dp_1 \LUT_reg[57][11]  ( .ip(n14389), .ck(clk), .q(\LUT[57][11] ) );
  dp_1 \LUT_reg[57][10]  ( .ip(n14388), .ck(clk), .q(\LUT[57][10] ) );
  dp_1 \LUT_reg[57][9]  ( .ip(n14387), .ck(clk), .q(\LUT[57][9] ) );
  dp_1 \LUT_reg[57][8]  ( .ip(n14386), .ck(clk), .q(\LUT[57][8] ) );
  dp_1 \LUT_reg[57][7]  ( .ip(n14385), .ck(clk), .q(\LUT[57][7] ) );
  dp_1 \LUT_reg[57][6]  ( .ip(n14384), .ck(clk), .q(\LUT[57][6] ) );
  dp_1 \LUT_reg[57][5]  ( .ip(n14383), .ck(clk), .q(\LUT[57][5] ) );
  dp_1 \LUT_reg[57][4]  ( .ip(n14382), .ck(clk), .q(\LUT[57][4] ) );
  dp_1 \LUT_reg[57][3]  ( .ip(n14381), .ck(clk), .q(\LUT[57][3] ) );
  dp_1 \LUT_reg[57][2]  ( .ip(n14380), .ck(clk), .q(\LUT[57][2] ) );
  dp_1 \LUT_reg[57][1]  ( .ip(n14379), .ck(clk), .q(\LUT[57][1] ) );
  dp_1 \LUT_reg[57][0]  ( .ip(n14378), .ck(clk), .q(\LUT[57][0] ) );
  dp_1 \LUT_reg[56][15]  ( .ip(n14377), .ck(clk), .q(\LUT[56][15] ) );
  dp_1 \LUT_reg[56][14]  ( .ip(n14376), .ck(clk), .q(\LUT[56][14] ) );
  dp_1 \LUT_reg[56][13]  ( .ip(n14375), .ck(clk), .q(\LUT[56][13] ) );
  dp_1 \LUT_reg[56][12]  ( .ip(n14374), .ck(clk), .q(\LUT[56][12] ) );
  dp_1 \LUT_reg[56][11]  ( .ip(n14373), .ck(clk), .q(\LUT[56][11] ) );
  dp_1 \LUT_reg[56][10]  ( .ip(n14372), .ck(clk), .q(\LUT[56][10] ) );
  dp_1 \LUT_reg[56][9]  ( .ip(n14371), .ck(clk), .q(\LUT[56][9] ) );
  dp_1 \LUT_reg[56][8]  ( .ip(n14370), .ck(clk), .q(\LUT[56][8] ) );
  dp_1 \LUT_reg[56][7]  ( .ip(n14369), .ck(clk), .q(\LUT[56][7] ) );
  dp_1 \LUT_reg[56][6]  ( .ip(n14368), .ck(clk), .q(\LUT[56][6] ) );
  dp_1 \LUT_reg[56][5]  ( .ip(n14367), .ck(clk), .q(\LUT[56][5] ) );
  dp_1 \LUT_reg[56][4]  ( .ip(n14366), .ck(clk), .q(\LUT[56][4] ) );
  dp_1 \LUT_reg[56][3]  ( .ip(n14365), .ck(clk), .q(\LUT[56][3] ) );
  dp_1 \LUT_reg[56][2]  ( .ip(n14364), .ck(clk), .q(\LUT[56][2] ) );
  dp_1 \LUT_reg[56][1]  ( .ip(n14363), .ck(clk), .q(\LUT[56][1] ) );
  dp_1 \LUT_reg[56][0]  ( .ip(n14362), .ck(clk), .q(\LUT[56][0] ) );
  dp_1 \LUT_reg[55][15]  ( .ip(n14361), .ck(clk), .q(\LUT[55][15] ) );
  dp_1 \LUT_reg[55][14]  ( .ip(n14360), .ck(clk), .q(\LUT[55][14] ) );
  dp_1 \LUT_reg[55][13]  ( .ip(n14359), .ck(clk), .q(\LUT[55][13] ) );
  dp_1 \LUT_reg[55][12]  ( .ip(n14358), .ck(clk), .q(\LUT[55][12] ) );
  dp_1 \LUT_reg[55][11]  ( .ip(n14357), .ck(clk), .q(\LUT[55][11] ) );
  dp_1 \LUT_reg[55][10]  ( .ip(n14356), .ck(clk), .q(\LUT[55][10] ) );
  dp_1 \LUT_reg[55][9]  ( .ip(n14355), .ck(clk), .q(\LUT[55][9] ) );
  dp_1 \LUT_reg[55][8]  ( .ip(n14354), .ck(clk), .q(\LUT[55][8] ) );
  dp_1 \LUT_reg[55][7]  ( .ip(n14353), .ck(clk), .q(\LUT[55][7] ) );
  dp_1 \LUT_reg[55][6]  ( .ip(n14352), .ck(clk), .q(\LUT[55][6] ) );
  dp_1 \LUT_reg[55][5]  ( .ip(n14351), .ck(clk), .q(\LUT[55][5] ) );
  dp_1 \LUT_reg[55][4]  ( .ip(n14350), .ck(clk), .q(\LUT[55][4] ) );
  dp_1 \LUT_reg[55][3]  ( .ip(n14349), .ck(clk), .q(\LUT[55][3] ) );
  dp_1 \LUT_reg[55][2]  ( .ip(n14348), .ck(clk), .q(\LUT[55][2] ) );
  dp_1 \LUT_reg[55][1]  ( .ip(n14347), .ck(clk), .q(\LUT[55][1] ) );
  dp_1 \LUT_reg[55][0]  ( .ip(n14346), .ck(clk), .q(\LUT[55][0] ) );
  dp_1 \LUT_reg[54][15]  ( .ip(n14345), .ck(clk), .q(\LUT[54][15] ) );
  dp_1 \LUT_reg[54][14]  ( .ip(n14344), .ck(clk), .q(\LUT[54][14] ) );
  dp_1 \LUT_reg[54][13]  ( .ip(n14343), .ck(clk), .q(\LUT[54][13] ) );
  dp_1 \LUT_reg[54][12]  ( .ip(n14342), .ck(clk), .q(\LUT[54][12] ) );
  dp_1 \LUT_reg[54][11]  ( .ip(n14341), .ck(clk), .q(\LUT[54][11] ) );
  dp_1 \LUT_reg[54][10]  ( .ip(n14340), .ck(clk), .q(\LUT[54][10] ) );
  dp_1 \LUT_reg[54][9]  ( .ip(n14339), .ck(clk), .q(\LUT[54][9] ) );
  dp_1 \LUT_reg[54][8]  ( .ip(n14338), .ck(clk), .q(\LUT[54][8] ) );
  dp_1 \LUT_reg[54][7]  ( .ip(n14337), .ck(clk), .q(\LUT[54][7] ) );
  dp_1 \LUT_reg[54][6]  ( .ip(n14336), .ck(clk), .q(\LUT[54][6] ) );
  dp_1 \LUT_reg[54][5]  ( .ip(n14335), .ck(clk), .q(\LUT[54][5] ) );
  dp_1 \LUT_reg[54][4]  ( .ip(n14334), .ck(clk), .q(\LUT[54][4] ) );
  dp_1 \LUT_reg[54][3]  ( .ip(n14333), .ck(clk), .q(\LUT[54][3] ) );
  dp_1 \LUT_reg[54][2]  ( .ip(n14332), .ck(clk), .q(\LUT[54][2] ) );
  dp_1 \LUT_reg[54][1]  ( .ip(n14331), .ck(clk), .q(\LUT[54][1] ) );
  dp_1 \LUT_reg[54][0]  ( .ip(n14330), .ck(clk), .q(\LUT[54][0] ) );
  dp_1 \LUT_reg[53][15]  ( .ip(n14329), .ck(clk), .q(\LUT[53][15] ) );
  dp_1 \LUT_reg[53][14]  ( .ip(n14328), .ck(clk), .q(\LUT[53][14] ) );
  dp_1 \LUT_reg[53][13]  ( .ip(n14327), .ck(clk), .q(\LUT[53][13] ) );
  dp_1 \LUT_reg[53][12]  ( .ip(n14326), .ck(clk), .q(\LUT[53][12] ) );
  dp_1 \LUT_reg[53][11]  ( .ip(n14325), .ck(clk), .q(\LUT[53][11] ) );
  dp_1 \LUT_reg[53][10]  ( .ip(n14324), .ck(clk), .q(\LUT[53][10] ) );
  dp_1 \LUT_reg[53][9]  ( .ip(n14323), .ck(clk), .q(\LUT[53][9] ) );
  dp_1 \LUT_reg[53][8]  ( .ip(n14322), .ck(clk), .q(\LUT[53][8] ) );
  dp_1 \LUT_reg[53][7]  ( .ip(n14321), .ck(clk), .q(\LUT[53][7] ) );
  dp_1 \LUT_reg[53][6]  ( .ip(n14320), .ck(clk), .q(\LUT[53][6] ) );
  dp_1 \LUT_reg[53][5]  ( .ip(n14319), .ck(clk), .q(\LUT[53][5] ) );
  dp_1 \LUT_reg[53][4]  ( .ip(n14318), .ck(clk), .q(\LUT[53][4] ) );
  dp_1 \LUT_reg[53][3]  ( .ip(n14317), .ck(clk), .q(\LUT[53][3] ) );
  dp_1 \LUT_reg[53][2]  ( .ip(n14316), .ck(clk), .q(\LUT[53][2] ) );
  dp_1 \LUT_reg[53][1]  ( .ip(n14315), .ck(clk), .q(\LUT[53][1] ) );
  dp_1 \LUT_reg[53][0]  ( .ip(n14314), .ck(clk), .q(\LUT[53][0] ) );
  dp_1 \LUT_reg[52][15]  ( .ip(n14313), .ck(clk), .q(\LUT[52][15] ) );
  dp_1 \LUT_reg[52][14]  ( .ip(n14312), .ck(clk), .q(\LUT[52][14] ) );
  dp_1 \LUT_reg[52][13]  ( .ip(n14311), .ck(clk), .q(\LUT[52][13] ) );
  dp_1 \LUT_reg[52][12]  ( .ip(n14310), .ck(clk), .q(\LUT[52][12] ) );
  dp_1 \LUT_reg[52][11]  ( .ip(n14309), .ck(clk), .q(\LUT[52][11] ) );
  dp_1 \LUT_reg[52][10]  ( .ip(n14308), .ck(clk), .q(\LUT[52][10] ) );
  dp_1 \LUT_reg[52][9]  ( .ip(n14307), .ck(clk), .q(\LUT[52][9] ) );
  dp_1 \LUT_reg[52][8]  ( .ip(n14306), .ck(clk), .q(\LUT[52][8] ) );
  dp_1 \LUT_reg[52][7]  ( .ip(n14305), .ck(clk), .q(\LUT[52][7] ) );
  dp_1 \LUT_reg[52][6]  ( .ip(n14304), .ck(clk), .q(\LUT[52][6] ) );
  dp_1 \LUT_reg[52][5]  ( .ip(n14303), .ck(clk), .q(\LUT[52][5] ) );
  dp_1 \LUT_reg[52][4]  ( .ip(n14302), .ck(clk), .q(\LUT[52][4] ) );
  dp_1 \LUT_reg[52][3]  ( .ip(n14301), .ck(clk), .q(\LUT[52][3] ) );
  dp_1 \LUT_reg[52][2]  ( .ip(n14300), .ck(clk), .q(\LUT[52][2] ) );
  dp_1 \LUT_reg[52][1]  ( .ip(n14299), .ck(clk), .q(\LUT[52][1] ) );
  dp_1 \LUT_reg[52][0]  ( .ip(n14298), .ck(clk), .q(\LUT[52][0] ) );
  dp_1 \LUT_reg[51][15]  ( .ip(n14297), .ck(clk), .q(\LUT[51][15] ) );
  dp_1 \LUT_reg[51][14]  ( .ip(n14296), .ck(clk), .q(\LUT[51][14] ) );
  dp_1 \LUT_reg[51][13]  ( .ip(n14295), .ck(clk), .q(\LUT[51][13] ) );
  dp_1 \LUT_reg[51][12]  ( .ip(n14294), .ck(clk), .q(\LUT[51][12] ) );
  dp_1 \LUT_reg[51][11]  ( .ip(n14293), .ck(clk), .q(\LUT[51][11] ) );
  dp_1 \LUT_reg[51][10]  ( .ip(n14292), .ck(clk), .q(\LUT[51][10] ) );
  dp_1 \LUT_reg[51][9]  ( .ip(n14291), .ck(clk), .q(\LUT[51][9] ) );
  dp_1 \LUT_reg[51][8]  ( .ip(n14290), .ck(clk), .q(\LUT[51][8] ) );
  dp_1 \LUT_reg[51][7]  ( .ip(n14289), .ck(clk), .q(\LUT[51][7] ) );
  dp_1 \LUT_reg[51][6]  ( .ip(n14288), .ck(clk), .q(\LUT[51][6] ) );
  dp_1 \LUT_reg[51][5]  ( .ip(n14287), .ck(clk), .q(\LUT[51][5] ) );
  dp_1 \LUT_reg[51][4]  ( .ip(n14286), .ck(clk), .q(\LUT[51][4] ) );
  dp_1 \LUT_reg[51][3]  ( .ip(n14285), .ck(clk), .q(\LUT[51][3] ) );
  dp_1 \LUT_reg[51][2]  ( .ip(n14284), .ck(clk), .q(\LUT[51][2] ) );
  dp_1 \LUT_reg[51][1]  ( .ip(n14283), .ck(clk), .q(\LUT[51][1] ) );
  dp_1 \LUT_reg[51][0]  ( .ip(n14282), .ck(clk), .q(\LUT[51][0] ) );
  dp_1 \LUT_reg[50][15]  ( .ip(n14281), .ck(clk), .q(\LUT[50][15] ) );
  dp_1 \LUT_reg[50][14]  ( .ip(n14280), .ck(clk), .q(\LUT[50][14] ) );
  dp_1 \LUT_reg[50][13]  ( .ip(n14279), .ck(clk), .q(\LUT[50][13] ) );
  dp_1 \LUT_reg[50][12]  ( .ip(n14278), .ck(clk), .q(\LUT[50][12] ) );
  dp_1 \LUT_reg[50][11]  ( .ip(n14277), .ck(clk), .q(\LUT[50][11] ) );
  dp_1 \LUT_reg[50][10]  ( .ip(n14276), .ck(clk), .q(\LUT[50][10] ) );
  dp_1 \LUT_reg[50][9]  ( .ip(n14275), .ck(clk), .q(\LUT[50][9] ) );
  dp_1 \LUT_reg[50][8]  ( .ip(n14274), .ck(clk), .q(\LUT[50][8] ) );
  dp_1 \LUT_reg[50][7]  ( .ip(n14273), .ck(clk), .q(\LUT[50][7] ) );
  dp_1 \LUT_reg[50][6]  ( .ip(n14272), .ck(clk), .q(\LUT[50][6] ) );
  dp_1 \LUT_reg[50][5]  ( .ip(n14271), .ck(clk), .q(\LUT[50][5] ) );
  dp_1 \LUT_reg[50][4]  ( .ip(n14270), .ck(clk), .q(\LUT[50][4] ) );
  dp_1 \LUT_reg[50][3]  ( .ip(n14269), .ck(clk), .q(\LUT[50][3] ) );
  dp_1 \LUT_reg[50][2]  ( .ip(n14268), .ck(clk), .q(\LUT[50][2] ) );
  dp_1 \LUT_reg[50][1]  ( .ip(n14267), .ck(clk), .q(\LUT[50][1] ) );
  dp_1 \LUT_reg[50][0]  ( .ip(n14266), .ck(clk), .q(\LUT[50][0] ) );
  dp_1 \LUT_reg[49][15]  ( .ip(n14265), .ck(clk), .q(\LUT[49][15] ) );
  dp_1 \LUT_reg[49][14]  ( .ip(n14264), .ck(clk), .q(\LUT[49][14] ) );
  dp_1 \LUT_reg[49][13]  ( .ip(n14263), .ck(clk), .q(\LUT[49][13] ) );
  dp_1 \LUT_reg[49][12]  ( .ip(n14262), .ck(clk), .q(\LUT[49][12] ) );
  dp_1 \LUT_reg[49][11]  ( .ip(n14261), .ck(clk), .q(\LUT[49][11] ) );
  dp_1 \LUT_reg[49][10]  ( .ip(n14260), .ck(clk), .q(\LUT[49][10] ) );
  dp_1 \LUT_reg[49][9]  ( .ip(n14259), .ck(clk), .q(\LUT[49][9] ) );
  dp_1 \LUT_reg[49][8]  ( .ip(n14258), .ck(clk), .q(\LUT[49][8] ) );
  dp_1 \LUT_reg[49][7]  ( .ip(n14257), .ck(clk), .q(\LUT[49][7] ) );
  dp_1 \LUT_reg[49][6]  ( .ip(n14256), .ck(clk), .q(\LUT[49][6] ) );
  dp_1 \LUT_reg[49][5]  ( .ip(n14255), .ck(clk), .q(\LUT[49][5] ) );
  dp_1 \LUT_reg[49][4]  ( .ip(n14254), .ck(clk), .q(\LUT[49][4] ) );
  dp_1 \LUT_reg[49][3]  ( .ip(n14253), .ck(clk), .q(\LUT[49][3] ) );
  dp_1 \LUT_reg[49][2]  ( .ip(n14252), .ck(clk), .q(\LUT[49][2] ) );
  dp_1 \LUT_reg[49][1]  ( .ip(n14251), .ck(clk), .q(\LUT[49][1] ) );
  dp_1 \LUT_reg[49][0]  ( .ip(n14250), .ck(clk), .q(\LUT[49][0] ) );
  dp_1 \LUT_reg[48][15]  ( .ip(n14249), .ck(clk), .q(\LUT[48][15] ) );
  dp_1 \LUT_reg[48][14]  ( .ip(n14248), .ck(clk), .q(\LUT[48][14] ) );
  dp_1 \LUT_reg[48][13]  ( .ip(n14247), .ck(clk), .q(\LUT[48][13] ) );
  dp_1 \LUT_reg[48][12]  ( .ip(n14246), .ck(clk), .q(\LUT[48][12] ) );
  dp_1 \LUT_reg[48][11]  ( .ip(n14245), .ck(clk), .q(\LUT[48][11] ) );
  dp_1 \LUT_reg[48][10]  ( .ip(n14244), .ck(clk), .q(\LUT[48][10] ) );
  dp_1 \LUT_reg[48][9]  ( .ip(n14243), .ck(clk), .q(\LUT[48][9] ) );
  dp_1 \LUT_reg[48][8]  ( .ip(n14242), .ck(clk), .q(\LUT[48][8] ) );
  dp_1 \LUT_reg[48][7]  ( .ip(n14241), .ck(clk), .q(\LUT[48][7] ) );
  dp_1 \LUT_reg[48][6]  ( .ip(n14240), .ck(clk), .q(\LUT[48][6] ) );
  dp_1 \LUT_reg[48][5]  ( .ip(n14239), .ck(clk), .q(\LUT[48][5] ) );
  dp_1 \LUT_reg[48][4]  ( .ip(n14238), .ck(clk), .q(\LUT[48][4] ) );
  dp_1 \LUT_reg[48][3]  ( .ip(n14237), .ck(clk), .q(\LUT[48][3] ) );
  dp_1 \LUT_reg[48][2]  ( .ip(n14236), .ck(clk), .q(\LUT[48][2] ) );
  dp_1 \LUT_reg[48][1]  ( .ip(n14235), .ck(clk), .q(\LUT[48][1] ) );
  dp_1 \LUT_reg[48][0]  ( .ip(n14234), .ck(clk), .q(\LUT[48][0] ) );
  dp_1 \LUT_reg[47][15]  ( .ip(n14233), .ck(clk), .q(\LUT[47][15] ) );
  dp_1 \LUT_reg[47][14]  ( .ip(n14232), .ck(clk), .q(\LUT[47][14] ) );
  dp_1 \LUT_reg[47][13]  ( .ip(n14231), .ck(clk), .q(\LUT[47][13] ) );
  dp_1 \LUT_reg[47][12]  ( .ip(n14230), .ck(clk), .q(\LUT[47][12] ) );
  dp_1 \LUT_reg[47][11]  ( .ip(n14229), .ck(clk), .q(\LUT[47][11] ) );
  dp_1 \LUT_reg[47][10]  ( .ip(n14228), .ck(clk), .q(\LUT[47][10] ) );
  dp_1 \LUT_reg[47][9]  ( .ip(n14227), .ck(clk), .q(\LUT[47][9] ) );
  dp_1 \LUT_reg[47][8]  ( .ip(n14226), .ck(clk), .q(\LUT[47][8] ) );
  dp_1 \LUT_reg[47][7]  ( .ip(n14225), .ck(clk), .q(\LUT[47][7] ) );
  dp_1 \LUT_reg[47][6]  ( .ip(n14224), .ck(clk), .q(\LUT[47][6] ) );
  dp_1 \LUT_reg[47][5]  ( .ip(n14223), .ck(clk), .q(\LUT[47][5] ) );
  dp_1 \LUT_reg[47][4]  ( .ip(n14222), .ck(clk), .q(\LUT[47][4] ) );
  dp_1 \LUT_reg[47][3]  ( .ip(n14221), .ck(clk), .q(\LUT[47][3] ) );
  dp_1 \LUT_reg[47][2]  ( .ip(n14220), .ck(clk), .q(\LUT[47][2] ) );
  dp_1 \LUT_reg[47][1]  ( .ip(n14219), .ck(clk), .q(\LUT[47][1] ) );
  dp_1 \LUT_reg[47][0]  ( .ip(n14218), .ck(clk), .q(\LUT[47][0] ) );
  dp_1 \LUT_reg[46][15]  ( .ip(n14217), .ck(clk), .q(\LUT[46][15] ) );
  dp_1 \LUT_reg[46][14]  ( .ip(n14216), .ck(clk), .q(\LUT[46][14] ) );
  dp_1 \LUT_reg[46][13]  ( .ip(n14215), .ck(clk), .q(\LUT[46][13] ) );
  dp_1 \LUT_reg[46][12]  ( .ip(n14214), .ck(clk), .q(\LUT[46][12] ) );
  dp_1 \LUT_reg[46][11]  ( .ip(n14213), .ck(clk), .q(\LUT[46][11] ) );
  dp_1 \LUT_reg[46][10]  ( .ip(n14212), .ck(clk), .q(\LUT[46][10] ) );
  dp_1 \LUT_reg[46][9]  ( .ip(n14211), .ck(clk), .q(\LUT[46][9] ) );
  dp_1 \LUT_reg[46][8]  ( .ip(n14210), .ck(clk), .q(\LUT[46][8] ) );
  dp_1 \LUT_reg[46][7]  ( .ip(n14209), .ck(clk), .q(\LUT[46][7] ) );
  dp_1 \LUT_reg[46][6]  ( .ip(n14208), .ck(clk), .q(\LUT[46][6] ) );
  dp_1 \LUT_reg[46][5]  ( .ip(n14207), .ck(clk), .q(\LUT[46][5] ) );
  dp_1 \LUT_reg[46][4]  ( .ip(n14206), .ck(clk), .q(\LUT[46][4] ) );
  dp_1 \LUT_reg[46][3]  ( .ip(n14205), .ck(clk), .q(\LUT[46][3] ) );
  dp_1 \LUT_reg[46][2]  ( .ip(n14204), .ck(clk), .q(\LUT[46][2] ) );
  dp_1 \LUT_reg[46][1]  ( .ip(n14203), .ck(clk), .q(\LUT[46][1] ) );
  dp_1 \LUT_reg[46][0]  ( .ip(n14202), .ck(clk), .q(\LUT[46][0] ) );
  dp_1 \LUT_reg[45][15]  ( .ip(n14201), .ck(clk), .q(\LUT[45][15] ) );
  dp_1 \LUT_reg[45][14]  ( .ip(n14200), .ck(clk), .q(\LUT[45][14] ) );
  dp_1 \LUT_reg[45][13]  ( .ip(n14199), .ck(clk), .q(\LUT[45][13] ) );
  dp_1 \LUT_reg[45][12]  ( .ip(n14198), .ck(clk), .q(\LUT[45][12] ) );
  dp_1 \LUT_reg[45][11]  ( .ip(n14197), .ck(clk), .q(\LUT[45][11] ) );
  dp_1 \LUT_reg[45][10]  ( .ip(n14196), .ck(clk), .q(\LUT[45][10] ) );
  dp_1 \LUT_reg[45][9]  ( .ip(n14195), .ck(clk), .q(\LUT[45][9] ) );
  dp_1 \LUT_reg[45][8]  ( .ip(n14194), .ck(clk), .q(\LUT[45][8] ) );
  dp_1 \LUT_reg[45][7]  ( .ip(n14193), .ck(clk), .q(\LUT[45][7] ) );
  dp_1 \LUT_reg[45][6]  ( .ip(n14192), .ck(clk), .q(\LUT[45][6] ) );
  dp_1 \LUT_reg[45][5]  ( .ip(n14191), .ck(clk), .q(\LUT[45][5] ) );
  dp_1 \LUT_reg[45][4]  ( .ip(n14190), .ck(clk), .q(\LUT[45][4] ) );
  dp_1 \LUT_reg[45][3]  ( .ip(n14189), .ck(clk), .q(\LUT[45][3] ) );
  dp_1 \LUT_reg[45][2]  ( .ip(n14188), .ck(clk), .q(\LUT[45][2] ) );
  dp_1 \LUT_reg[45][1]  ( .ip(n14187), .ck(clk), .q(\LUT[45][1] ) );
  dp_1 \LUT_reg[45][0]  ( .ip(n14186), .ck(clk), .q(\LUT[45][0] ) );
  dp_1 \LUT_reg[44][15]  ( .ip(n14185), .ck(clk), .q(\LUT[44][15] ) );
  dp_1 \LUT_reg[44][14]  ( .ip(n14184), .ck(clk), .q(\LUT[44][14] ) );
  dp_1 \LUT_reg[44][13]  ( .ip(n14183), .ck(clk), .q(\LUT[44][13] ) );
  dp_1 \LUT_reg[44][12]  ( .ip(n14182), .ck(clk), .q(\LUT[44][12] ) );
  dp_1 \LUT_reg[44][11]  ( .ip(n14181), .ck(clk), .q(\LUT[44][11] ) );
  dp_1 \LUT_reg[44][10]  ( .ip(n14180), .ck(clk), .q(\LUT[44][10] ) );
  dp_1 \LUT_reg[44][9]  ( .ip(n14179), .ck(clk), .q(\LUT[44][9] ) );
  dp_1 \LUT_reg[44][8]  ( .ip(n14178), .ck(clk), .q(\LUT[44][8] ) );
  dp_1 \LUT_reg[44][7]  ( .ip(n14177), .ck(clk), .q(\LUT[44][7] ) );
  dp_1 \LUT_reg[44][6]  ( .ip(n14176), .ck(clk), .q(\LUT[44][6] ) );
  dp_1 \LUT_reg[44][5]  ( .ip(n14175), .ck(clk), .q(\LUT[44][5] ) );
  dp_1 \LUT_reg[44][4]  ( .ip(n14174), .ck(clk), .q(\LUT[44][4] ) );
  dp_1 \LUT_reg[44][3]  ( .ip(n14173), .ck(clk), .q(\LUT[44][3] ) );
  dp_1 \LUT_reg[44][2]  ( .ip(n14172), .ck(clk), .q(\LUT[44][2] ) );
  dp_1 \LUT_reg[44][1]  ( .ip(n14171), .ck(clk), .q(\LUT[44][1] ) );
  dp_1 \LUT_reg[44][0]  ( .ip(n14170), .ck(clk), .q(\LUT[44][0] ) );
  dp_1 \LUT_reg[43][15]  ( .ip(n14169), .ck(clk), .q(\LUT[43][15] ) );
  dp_1 \LUT_reg[43][14]  ( .ip(n14168), .ck(clk), .q(\LUT[43][14] ) );
  dp_1 \LUT_reg[43][13]  ( .ip(n14167), .ck(clk), .q(\LUT[43][13] ) );
  dp_1 \LUT_reg[43][12]  ( .ip(n14166), .ck(clk), .q(\LUT[43][12] ) );
  dp_1 \LUT_reg[43][11]  ( .ip(n14165), .ck(clk), .q(\LUT[43][11] ) );
  dp_1 \LUT_reg[43][10]  ( .ip(n14164), .ck(clk), .q(\LUT[43][10] ) );
  dp_1 \LUT_reg[43][9]  ( .ip(n14163), .ck(clk), .q(\LUT[43][9] ) );
  dp_1 \LUT_reg[43][8]  ( .ip(n14162), .ck(clk), .q(\LUT[43][8] ) );
  dp_1 \LUT_reg[43][7]  ( .ip(n14161), .ck(clk), .q(\LUT[43][7] ) );
  dp_1 \LUT_reg[43][6]  ( .ip(n14160), .ck(clk), .q(\LUT[43][6] ) );
  dp_1 \LUT_reg[43][5]  ( .ip(n14159), .ck(clk), .q(\LUT[43][5] ) );
  dp_1 \LUT_reg[43][4]  ( .ip(n14158), .ck(clk), .q(\LUT[43][4] ) );
  dp_1 \LUT_reg[43][3]  ( .ip(n14157), .ck(clk), .q(\LUT[43][3] ) );
  dp_1 \LUT_reg[43][2]  ( .ip(n14156), .ck(clk), .q(\LUT[43][2] ) );
  dp_1 \LUT_reg[43][1]  ( .ip(n14155), .ck(clk), .q(\LUT[43][1] ) );
  dp_1 \LUT_reg[43][0]  ( .ip(n14154), .ck(clk), .q(\LUT[43][0] ) );
  dp_1 \LUT_reg[42][15]  ( .ip(n14153), .ck(clk), .q(\LUT[42][15] ) );
  dp_1 \LUT_reg[42][14]  ( .ip(n14152), .ck(clk), .q(\LUT[42][14] ) );
  dp_1 \LUT_reg[42][13]  ( .ip(n14151), .ck(clk), .q(\LUT[42][13] ) );
  dp_1 \LUT_reg[42][12]  ( .ip(n14150), .ck(clk), .q(\LUT[42][12] ) );
  dp_1 \LUT_reg[42][11]  ( .ip(n14149), .ck(clk), .q(\LUT[42][11] ) );
  dp_1 \LUT_reg[42][10]  ( .ip(n14148), .ck(clk), .q(\LUT[42][10] ) );
  dp_1 \LUT_reg[42][9]  ( .ip(n14147), .ck(clk), .q(\LUT[42][9] ) );
  dp_1 \LUT_reg[42][8]  ( .ip(n14146), .ck(clk), .q(\LUT[42][8] ) );
  dp_1 \LUT_reg[42][7]  ( .ip(n14145), .ck(clk), .q(\LUT[42][7] ) );
  dp_1 \LUT_reg[42][6]  ( .ip(n14144), .ck(clk), .q(\LUT[42][6] ) );
  dp_1 \LUT_reg[42][5]  ( .ip(n14143), .ck(clk), .q(\LUT[42][5] ) );
  dp_1 \LUT_reg[42][4]  ( .ip(n14142), .ck(clk), .q(\LUT[42][4] ) );
  dp_1 \LUT_reg[42][3]  ( .ip(n14141), .ck(clk), .q(\LUT[42][3] ) );
  dp_1 \LUT_reg[42][2]  ( .ip(n14140), .ck(clk), .q(\LUT[42][2] ) );
  dp_1 \LUT_reg[42][1]  ( .ip(n14139), .ck(clk), .q(\LUT[42][1] ) );
  dp_1 \LUT_reg[42][0]  ( .ip(n14138), .ck(clk), .q(\LUT[42][0] ) );
  dp_1 \LUT_reg[41][15]  ( .ip(n14137), .ck(clk), .q(\LUT[41][15] ) );
  dp_1 \LUT_reg[41][14]  ( .ip(n14136), .ck(clk), .q(\LUT[41][14] ) );
  dp_1 \LUT_reg[41][13]  ( .ip(n14135), .ck(clk), .q(\LUT[41][13] ) );
  dp_1 \LUT_reg[41][12]  ( .ip(n14134), .ck(clk), .q(\LUT[41][12] ) );
  dp_1 \LUT_reg[41][11]  ( .ip(n14133), .ck(clk), .q(\LUT[41][11] ) );
  dp_1 \LUT_reg[41][10]  ( .ip(n14132), .ck(clk), .q(\LUT[41][10] ) );
  dp_1 \LUT_reg[41][9]  ( .ip(n14131), .ck(clk), .q(\LUT[41][9] ) );
  dp_1 \LUT_reg[41][8]  ( .ip(n14130), .ck(clk), .q(\LUT[41][8] ) );
  dp_1 \LUT_reg[41][7]  ( .ip(n14129), .ck(clk), .q(\LUT[41][7] ) );
  dp_1 \LUT_reg[41][6]  ( .ip(n14128), .ck(clk), .q(\LUT[41][6] ) );
  dp_1 \LUT_reg[41][5]  ( .ip(n14127), .ck(clk), .q(\LUT[41][5] ) );
  dp_1 \LUT_reg[41][4]  ( .ip(n14126), .ck(clk), .q(\LUT[41][4] ) );
  dp_1 \LUT_reg[41][3]  ( .ip(n14125), .ck(clk), .q(\LUT[41][3] ) );
  dp_1 \LUT_reg[41][2]  ( .ip(n14124), .ck(clk), .q(\LUT[41][2] ) );
  dp_1 \LUT_reg[41][1]  ( .ip(n14123), .ck(clk), .q(\LUT[41][1] ) );
  dp_1 \LUT_reg[41][0]  ( .ip(n14122), .ck(clk), .q(\LUT[41][0] ) );
  dp_1 \LUT_reg[40][15]  ( .ip(n14121), .ck(clk), .q(\LUT[40][15] ) );
  dp_1 \LUT_reg[40][14]  ( .ip(n14120), .ck(clk), .q(\LUT[40][14] ) );
  dp_1 \LUT_reg[40][13]  ( .ip(n14119), .ck(clk), .q(\LUT[40][13] ) );
  dp_1 \LUT_reg[40][12]  ( .ip(n14118), .ck(clk), .q(\LUT[40][12] ) );
  dp_1 \LUT_reg[40][11]  ( .ip(n14117), .ck(clk), .q(\LUT[40][11] ) );
  dp_1 \LUT_reg[40][10]  ( .ip(n14116), .ck(clk), .q(\LUT[40][10] ) );
  dp_1 \LUT_reg[40][9]  ( .ip(n14115), .ck(clk), .q(\LUT[40][9] ) );
  dp_1 \LUT_reg[40][8]  ( .ip(n14114), .ck(clk), .q(\LUT[40][8] ) );
  dp_1 \LUT_reg[40][7]  ( .ip(n14113), .ck(clk), .q(\LUT[40][7] ) );
  dp_1 \LUT_reg[40][6]  ( .ip(n14112), .ck(clk), .q(\LUT[40][6] ) );
  dp_1 \LUT_reg[40][5]  ( .ip(n14111), .ck(clk), .q(\LUT[40][5] ) );
  dp_1 \LUT_reg[40][4]  ( .ip(n14110), .ck(clk), .q(\LUT[40][4] ) );
  dp_1 \LUT_reg[40][3]  ( .ip(n14109), .ck(clk), .q(\LUT[40][3] ) );
  dp_1 \LUT_reg[40][2]  ( .ip(n14108), .ck(clk), .q(\LUT[40][2] ) );
  dp_1 \LUT_reg[40][1]  ( .ip(n14107), .ck(clk), .q(\LUT[40][1] ) );
  dp_1 \LUT_reg[40][0]  ( .ip(n14106), .ck(clk), .q(\LUT[40][0] ) );
  dp_1 \LUT_reg[39][15]  ( .ip(n14105), .ck(clk), .q(\LUT[39][15] ) );
  dp_1 \LUT_reg[39][14]  ( .ip(n14104), .ck(clk), .q(\LUT[39][14] ) );
  dp_1 \LUT_reg[39][13]  ( .ip(n14103), .ck(clk), .q(\LUT[39][13] ) );
  dp_1 \LUT_reg[39][12]  ( .ip(n14102), .ck(clk), .q(\LUT[39][12] ) );
  dp_1 \LUT_reg[39][11]  ( .ip(n14101), .ck(clk), .q(\LUT[39][11] ) );
  dp_1 \LUT_reg[39][10]  ( .ip(n14100), .ck(clk), .q(\LUT[39][10] ) );
  dp_1 \LUT_reg[39][9]  ( .ip(n14099), .ck(clk), .q(\LUT[39][9] ) );
  dp_1 \LUT_reg[39][8]  ( .ip(n14098), .ck(clk), .q(\LUT[39][8] ) );
  dp_1 \LUT_reg[39][7]  ( .ip(n14097), .ck(clk), .q(\LUT[39][7] ) );
  dp_1 \LUT_reg[39][6]  ( .ip(n14096), .ck(clk), .q(\LUT[39][6] ) );
  dp_1 \LUT_reg[39][5]  ( .ip(n14095), .ck(clk), .q(\LUT[39][5] ) );
  dp_1 \LUT_reg[39][4]  ( .ip(n14094), .ck(clk), .q(\LUT[39][4] ) );
  dp_1 \LUT_reg[39][3]  ( .ip(n14093), .ck(clk), .q(\LUT[39][3] ) );
  dp_1 \LUT_reg[39][2]  ( .ip(n14092), .ck(clk), .q(\LUT[39][2] ) );
  dp_1 \LUT_reg[39][1]  ( .ip(n14091), .ck(clk), .q(\LUT[39][1] ) );
  dp_1 \LUT_reg[39][0]  ( .ip(n14090), .ck(clk), .q(\LUT[39][0] ) );
  dp_1 \LUT_reg[38][15]  ( .ip(n14089), .ck(clk), .q(\LUT[38][15] ) );
  dp_1 \LUT_reg[38][14]  ( .ip(n14088), .ck(clk), .q(\LUT[38][14] ) );
  dp_1 \LUT_reg[38][13]  ( .ip(n14087), .ck(clk), .q(\LUT[38][13] ) );
  dp_1 \LUT_reg[38][12]  ( .ip(n14086), .ck(clk), .q(\LUT[38][12] ) );
  dp_1 \LUT_reg[38][11]  ( .ip(n14085), .ck(clk), .q(\LUT[38][11] ) );
  dp_1 \LUT_reg[38][10]  ( .ip(n14084), .ck(clk), .q(\LUT[38][10] ) );
  dp_1 \LUT_reg[38][9]  ( .ip(n14083), .ck(clk), .q(\LUT[38][9] ) );
  dp_1 \LUT_reg[38][8]  ( .ip(n14082), .ck(clk), .q(\LUT[38][8] ) );
  dp_1 \LUT_reg[38][7]  ( .ip(n14081), .ck(clk), .q(\LUT[38][7] ) );
  dp_1 \LUT_reg[38][6]  ( .ip(n14080), .ck(clk), .q(\LUT[38][6] ) );
  dp_1 \LUT_reg[38][5]  ( .ip(n14079), .ck(clk), .q(\LUT[38][5] ) );
  dp_1 \LUT_reg[38][4]  ( .ip(n14078), .ck(clk), .q(\LUT[38][4] ) );
  dp_1 \LUT_reg[38][3]  ( .ip(n14077), .ck(clk), .q(\LUT[38][3] ) );
  dp_1 \LUT_reg[38][2]  ( .ip(n14076), .ck(clk), .q(\LUT[38][2] ) );
  dp_1 \LUT_reg[38][1]  ( .ip(n14075), .ck(clk), .q(\LUT[38][1] ) );
  dp_1 \LUT_reg[38][0]  ( .ip(n14074), .ck(clk), .q(\LUT[38][0] ) );
  dp_1 \LUT_reg[37][15]  ( .ip(n14073), .ck(clk), .q(\LUT[37][15] ) );
  dp_1 \LUT_reg[37][14]  ( .ip(n14072), .ck(clk), .q(\LUT[37][14] ) );
  dp_1 \LUT_reg[37][13]  ( .ip(n14071), .ck(clk), .q(\LUT[37][13] ) );
  dp_1 \LUT_reg[37][12]  ( .ip(n14070), .ck(clk), .q(\LUT[37][12] ) );
  dp_1 \LUT_reg[37][11]  ( .ip(n14069), .ck(clk), .q(\LUT[37][11] ) );
  dp_1 \LUT_reg[37][10]  ( .ip(n14068), .ck(clk), .q(\LUT[37][10] ) );
  dp_1 \LUT_reg[37][9]  ( .ip(n14067), .ck(clk), .q(\LUT[37][9] ) );
  dp_1 \LUT_reg[37][8]  ( .ip(n14066), .ck(clk), .q(\LUT[37][8] ) );
  dp_1 \LUT_reg[37][7]  ( .ip(n14065), .ck(clk), .q(\LUT[37][7] ) );
  dp_1 \LUT_reg[37][6]  ( .ip(n14064), .ck(clk), .q(\LUT[37][6] ) );
  dp_1 \LUT_reg[37][5]  ( .ip(n14063), .ck(clk), .q(\LUT[37][5] ) );
  dp_1 \LUT_reg[37][4]  ( .ip(n14062), .ck(clk), .q(\LUT[37][4] ) );
  dp_1 \LUT_reg[37][3]  ( .ip(n14061), .ck(clk), .q(\LUT[37][3] ) );
  dp_1 \LUT_reg[37][2]  ( .ip(n14060), .ck(clk), .q(\LUT[37][2] ) );
  dp_1 \LUT_reg[37][1]  ( .ip(n14059), .ck(clk), .q(\LUT[37][1] ) );
  dp_1 \LUT_reg[37][0]  ( .ip(n14058), .ck(clk), .q(\LUT[37][0] ) );
  dp_1 \LUT_reg[36][15]  ( .ip(n14057), .ck(clk), .q(\LUT[36][15] ) );
  dp_1 \LUT_reg[36][14]  ( .ip(n14056), .ck(clk), .q(\LUT[36][14] ) );
  dp_1 \LUT_reg[36][13]  ( .ip(n14055), .ck(clk), .q(\LUT[36][13] ) );
  dp_1 \LUT_reg[36][12]  ( .ip(n14054), .ck(clk), .q(\LUT[36][12] ) );
  dp_1 \LUT_reg[36][11]  ( .ip(n14053), .ck(clk), .q(\LUT[36][11] ) );
  dp_1 \LUT_reg[36][10]  ( .ip(n14052), .ck(clk), .q(\LUT[36][10] ) );
  dp_1 \LUT_reg[36][9]  ( .ip(n14051), .ck(clk), .q(\LUT[36][9] ) );
  dp_1 \LUT_reg[36][8]  ( .ip(n14050), .ck(clk), .q(\LUT[36][8] ) );
  dp_1 \LUT_reg[36][7]  ( .ip(n14049), .ck(clk), .q(\LUT[36][7] ) );
  dp_1 \LUT_reg[36][6]  ( .ip(n14048), .ck(clk), .q(\LUT[36][6] ) );
  dp_1 \LUT_reg[36][5]  ( .ip(n14047), .ck(clk), .q(\LUT[36][5] ) );
  dp_1 \LUT_reg[36][4]  ( .ip(n14046), .ck(clk), .q(\LUT[36][4] ) );
  dp_1 \LUT_reg[36][3]  ( .ip(n14045), .ck(clk), .q(\LUT[36][3] ) );
  dp_1 \LUT_reg[36][2]  ( .ip(n14044), .ck(clk), .q(\LUT[36][2] ) );
  dp_1 \LUT_reg[36][1]  ( .ip(n14043), .ck(clk), .q(\LUT[36][1] ) );
  dp_1 \LUT_reg[36][0]  ( .ip(n14042), .ck(clk), .q(\LUT[36][0] ) );
  dp_1 \LUT_reg[35][15]  ( .ip(n14041), .ck(clk), .q(\LUT[35][15] ) );
  dp_1 \LUT_reg[35][14]  ( .ip(n14040), .ck(clk), .q(\LUT[35][14] ) );
  dp_1 \LUT_reg[35][13]  ( .ip(n14039), .ck(clk), .q(\LUT[35][13] ) );
  dp_1 \LUT_reg[35][12]  ( .ip(n14038), .ck(clk), .q(\LUT[35][12] ) );
  dp_1 \LUT_reg[35][11]  ( .ip(n14037), .ck(clk), .q(\LUT[35][11] ) );
  dp_1 \LUT_reg[35][10]  ( .ip(n14036), .ck(clk), .q(\LUT[35][10] ) );
  dp_1 \LUT_reg[35][9]  ( .ip(n14035), .ck(clk), .q(\LUT[35][9] ) );
  dp_1 \LUT_reg[35][8]  ( .ip(n14034), .ck(clk), .q(\LUT[35][8] ) );
  dp_1 \LUT_reg[35][7]  ( .ip(n14033), .ck(clk), .q(\LUT[35][7] ) );
  dp_1 \LUT_reg[35][6]  ( .ip(n14032), .ck(clk), .q(\LUT[35][6] ) );
  dp_1 \LUT_reg[35][5]  ( .ip(n14031), .ck(clk), .q(\LUT[35][5] ) );
  dp_1 \LUT_reg[35][4]  ( .ip(n14030), .ck(clk), .q(\LUT[35][4] ) );
  dp_1 \LUT_reg[35][3]  ( .ip(n14029), .ck(clk), .q(\LUT[35][3] ) );
  dp_1 \LUT_reg[35][2]  ( .ip(n14028), .ck(clk), .q(\LUT[35][2] ) );
  dp_1 \LUT_reg[35][1]  ( .ip(n14027), .ck(clk), .q(\LUT[35][1] ) );
  dp_1 \LUT_reg[35][0]  ( .ip(n14026), .ck(clk), .q(\LUT[35][0] ) );
  dp_1 \LUT_reg[34][15]  ( .ip(n14025), .ck(clk), .q(\LUT[34][15] ) );
  dp_1 \LUT_reg[34][14]  ( .ip(n14024), .ck(clk), .q(\LUT[34][14] ) );
  dp_1 \LUT_reg[34][13]  ( .ip(n14023), .ck(clk), .q(\LUT[34][13] ) );
  dp_1 \LUT_reg[34][12]  ( .ip(n14022), .ck(clk), .q(\LUT[34][12] ) );
  dp_1 \LUT_reg[34][11]  ( .ip(n14021), .ck(clk), .q(\LUT[34][11] ) );
  dp_1 \LUT_reg[34][10]  ( .ip(n14020), .ck(clk), .q(\LUT[34][10] ) );
  dp_1 \LUT_reg[34][9]  ( .ip(n14019), .ck(clk), .q(\LUT[34][9] ) );
  dp_1 \LUT_reg[34][8]  ( .ip(n14018), .ck(clk), .q(\LUT[34][8] ) );
  dp_1 \LUT_reg[34][7]  ( .ip(n14017), .ck(clk), .q(\LUT[34][7] ) );
  dp_1 \LUT_reg[34][6]  ( .ip(n14016), .ck(clk), .q(\LUT[34][6] ) );
  dp_1 \LUT_reg[34][5]  ( .ip(n14015), .ck(clk), .q(\LUT[34][5] ) );
  dp_1 \LUT_reg[34][4]  ( .ip(n14014), .ck(clk), .q(\LUT[34][4] ) );
  dp_1 \LUT_reg[34][3]  ( .ip(n14013), .ck(clk), .q(\LUT[34][3] ) );
  dp_1 \LUT_reg[34][2]  ( .ip(n14012), .ck(clk), .q(\LUT[34][2] ) );
  dp_1 \LUT_reg[34][1]  ( .ip(n14011), .ck(clk), .q(\LUT[34][1] ) );
  dp_1 \LUT_reg[34][0]  ( .ip(n14010), .ck(clk), .q(\LUT[34][0] ) );
  dp_1 \LUT_reg[33][15]  ( .ip(n14009), .ck(clk), .q(\LUT[33][15] ) );
  dp_1 \LUT_reg[33][14]  ( .ip(n14008), .ck(clk), .q(\LUT[33][14] ) );
  dp_1 \LUT_reg[33][13]  ( .ip(n14007), .ck(clk), .q(\LUT[33][13] ) );
  dp_1 \LUT_reg[33][12]  ( .ip(n14006), .ck(clk), .q(\LUT[33][12] ) );
  dp_1 \LUT_reg[33][11]  ( .ip(n14005), .ck(clk), .q(\LUT[33][11] ) );
  dp_1 \LUT_reg[33][10]  ( .ip(n14004), .ck(clk), .q(\LUT[33][10] ) );
  dp_1 \LUT_reg[33][9]  ( .ip(n14003), .ck(clk), .q(\LUT[33][9] ) );
  dp_1 \LUT_reg[33][8]  ( .ip(n14002), .ck(clk), .q(\LUT[33][8] ) );
  dp_1 \LUT_reg[33][7]  ( .ip(n14001), .ck(clk), .q(\LUT[33][7] ) );
  dp_1 \LUT_reg[33][6]  ( .ip(n14000), .ck(clk), .q(\LUT[33][6] ) );
  dp_1 \LUT_reg[33][5]  ( .ip(n13999), .ck(clk), .q(\LUT[33][5] ) );
  dp_1 \LUT_reg[33][4]  ( .ip(n13998), .ck(clk), .q(\LUT[33][4] ) );
  dp_1 \LUT_reg[33][3]  ( .ip(n13997), .ck(clk), .q(\LUT[33][3] ) );
  dp_1 \LUT_reg[33][2]  ( .ip(n13996), .ck(clk), .q(\LUT[33][2] ) );
  dp_1 \LUT_reg[33][1]  ( .ip(n13995), .ck(clk), .q(\LUT[33][1] ) );
  dp_1 \LUT_reg[33][0]  ( .ip(n13994), .ck(clk), .q(\LUT[33][0] ) );
  dp_1 \LUT_reg[32][15]  ( .ip(n13993), .ck(clk), .q(\LUT[32][15] ) );
  dp_1 \LUT_reg[32][14]  ( .ip(n13992), .ck(clk), .q(\LUT[32][14] ) );
  dp_1 \LUT_reg[32][13]  ( .ip(n13991), .ck(clk), .q(\LUT[32][13] ) );
  dp_1 \LUT_reg[32][12]  ( .ip(n13990), .ck(clk), .q(\LUT[32][12] ) );
  dp_1 \LUT_reg[32][11]  ( .ip(n13989), .ck(clk), .q(\LUT[32][11] ) );
  dp_1 \LUT_reg[32][10]  ( .ip(n13988), .ck(clk), .q(\LUT[32][10] ) );
  dp_1 \LUT_reg[32][9]  ( .ip(n13987), .ck(clk), .q(\LUT[32][9] ) );
  dp_1 \LUT_reg[32][8]  ( .ip(n13986), .ck(clk), .q(\LUT[32][8] ) );
  dp_1 \LUT_reg[32][7]  ( .ip(n13985), .ck(clk), .q(\LUT[32][7] ) );
  dp_1 \LUT_reg[32][6]  ( .ip(n13984), .ck(clk), .q(\LUT[32][6] ) );
  dp_1 \LUT_reg[32][5]  ( .ip(n13983), .ck(clk), .q(\LUT[32][5] ) );
  dp_1 \LUT_reg[32][4]  ( .ip(n13982), .ck(clk), .q(\LUT[32][4] ) );
  dp_1 \LUT_reg[32][3]  ( .ip(n13981), .ck(clk), .q(\LUT[32][3] ) );
  dp_1 \LUT_reg[32][2]  ( .ip(n13980), .ck(clk), .q(\LUT[32][2] ) );
  dp_1 \LUT_reg[32][1]  ( .ip(n13979), .ck(clk), .q(\LUT[32][1] ) );
  dp_1 \LUT_reg[32][0]  ( .ip(n13978), .ck(clk), .q(\LUT[32][0] ) );
  dp_1 \LUT_reg[31][15]  ( .ip(n13977), .ck(clk), .q(\LUT[31][15] ) );
  dp_1 \LUT_reg[31][14]  ( .ip(n13976), .ck(clk), .q(\LUT[31][14] ) );
  dp_1 \LUT_reg[31][13]  ( .ip(n13975), .ck(clk), .q(\LUT[31][13] ) );
  dp_1 \LUT_reg[31][12]  ( .ip(n13974), .ck(clk), .q(\LUT[31][12] ) );
  dp_1 \LUT_reg[31][11]  ( .ip(n13973), .ck(clk), .q(\LUT[31][11] ) );
  dp_1 \LUT_reg[31][10]  ( .ip(n13972), .ck(clk), .q(\LUT[31][10] ) );
  dp_1 \LUT_reg[31][9]  ( .ip(n13971), .ck(clk), .q(\LUT[31][9] ) );
  dp_1 \LUT_reg[31][8]  ( .ip(n13970), .ck(clk), .q(\LUT[31][8] ) );
  dp_1 \LUT_reg[31][7]  ( .ip(n13969), .ck(clk), .q(\LUT[31][7] ) );
  dp_1 \LUT_reg[31][6]  ( .ip(n13968), .ck(clk), .q(\LUT[31][6] ) );
  dp_1 \LUT_reg[31][5]  ( .ip(n13967), .ck(clk), .q(\LUT[31][5] ) );
  dp_1 \LUT_reg[31][4]  ( .ip(n13966), .ck(clk), .q(\LUT[31][4] ) );
  dp_1 \LUT_reg[31][3]  ( .ip(n13965), .ck(clk), .q(\LUT[31][3] ) );
  dp_1 \LUT_reg[31][2]  ( .ip(n13964), .ck(clk), .q(\LUT[31][2] ) );
  dp_1 \LUT_reg[31][1]  ( .ip(n13963), .ck(clk), .q(\LUT[31][1] ) );
  dp_1 \LUT_reg[31][0]  ( .ip(n13962), .ck(clk), .q(\LUT[31][0] ) );
  dp_1 \LUT_reg[30][15]  ( .ip(n13961), .ck(clk), .q(\LUT[30][15] ) );
  dp_1 \LUT_reg[30][14]  ( .ip(n13960), .ck(clk), .q(\LUT[30][14] ) );
  dp_1 \LUT_reg[30][13]  ( .ip(n13959), .ck(clk), .q(\LUT[30][13] ) );
  dp_1 \LUT_reg[30][12]  ( .ip(n13958), .ck(clk), .q(\LUT[30][12] ) );
  dp_1 \LUT_reg[30][11]  ( .ip(n13957), .ck(clk), .q(\LUT[30][11] ) );
  dp_1 \LUT_reg[30][10]  ( .ip(n13956), .ck(clk), .q(\LUT[30][10] ) );
  dp_1 \LUT_reg[30][9]  ( .ip(n13955), .ck(clk), .q(\LUT[30][9] ) );
  dp_1 \LUT_reg[30][8]  ( .ip(n13954), .ck(clk), .q(\LUT[30][8] ) );
  dp_1 \LUT_reg[30][7]  ( .ip(n13953), .ck(clk), .q(\LUT[30][7] ) );
  dp_1 \LUT_reg[30][6]  ( .ip(n13952), .ck(clk), .q(\LUT[30][6] ) );
  dp_1 \LUT_reg[30][5]  ( .ip(n13951), .ck(clk), .q(\LUT[30][5] ) );
  dp_1 \LUT_reg[30][4]  ( .ip(n13950), .ck(clk), .q(\LUT[30][4] ) );
  dp_1 \LUT_reg[30][3]  ( .ip(n13949), .ck(clk), .q(\LUT[30][3] ) );
  dp_1 \LUT_reg[30][2]  ( .ip(n13948), .ck(clk), .q(\LUT[30][2] ) );
  dp_1 \LUT_reg[30][1]  ( .ip(n13947), .ck(clk), .q(\LUT[30][1] ) );
  dp_1 \LUT_reg[30][0]  ( .ip(n13946), .ck(clk), .q(\LUT[30][0] ) );
  dp_1 \LUT_reg[29][15]  ( .ip(n13945), .ck(clk), .q(\LUT[29][15] ) );
  dp_1 \LUT_reg[29][14]  ( .ip(n13944), .ck(clk), .q(\LUT[29][14] ) );
  dp_1 \LUT_reg[29][13]  ( .ip(n13943), .ck(clk), .q(\LUT[29][13] ) );
  dp_1 \LUT_reg[29][12]  ( .ip(n13942), .ck(clk), .q(\LUT[29][12] ) );
  dp_1 \LUT_reg[29][11]  ( .ip(n13941), .ck(clk), .q(\LUT[29][11] ) );
  dp_1 \LUT_reg[29][10]  ( .ip(n13940), .ck(clk), .q(\LUT[29][10] ) );
  dp_1 \LUT_reg[29][9]  ( .ip(n13939), .ck(clk), .q(\LUT[29][9] ) );
  dp_1 \LUT_reg[29][8]  ( .ip(n13938), .ck(clk), .q(\LUT[29][8] ) );
  dp_1 \LUT_reg[29][7]  ( .ip(n13937), .ck(clk), .q(\LUT[29][7] ) );
  dp_1 \LUT_reg[29][6]  ( .ip(n13936), .ck(clk), .q(\LUT[29][6] ) );
  dp_1 \LUT_reg[29][5]  ( .ip(n13935), .ck(clk), .q(\LUT[29][5] ) );
  dp_1 \LUT_reg[29][4]  ( .ip(n13934), .ck(clk), .q(\LUT[29][4] ) );
  dp_1 \LUT_reg[29][3]  ( .ip(n13933), .ck(clk), .q(\LUT[29][3] ) );
  dp_1 \LUT_reg[29][2]  ( .ip(n13932), .ck(clk), .q(\LUT[29][2] ) );
  dp_1 \LUT_reg[29][1]  ( .ip(n13931), .ck(clk), .q(\LUT[29][1] ) );
  dp_1 \LUT_reg[29][0]  ( .ip(n13930), .ck(clk), .q(\LUT[29][0] ) );
  dp_1 \LUT_reg[28][15]  ( .ip(n13929), .ck(clk), .q(\LUT[28][15] ) );
  dp_1 \LUT_reg[28][14]  ( .ip(n13928), .ck(clk), .q(\LUT[28][14] ) );
  dp_1 \LUT_reg[28][13]  ( .ip(n13927), .ck(clk), .q(\LUT[28][13] ) );
  dp_1 \LUT_reg[28][12]  ( .ip(n13926), .ck(clk), .q(\LUT[28][12] ) );
  dp_1 \LUT_reg[28][11]  ( .ip(n13925), .ck(clk), .q(\LUT[28][11] ) );
  dp_1 \LUT_reg[28][10]  ( .ip(n13924), .ck(clk), .q(\LUT[28][10] ) );
  dp_1 \LUT_reg[28][9]  ( .ip(n13923), .ck(clk), .q(\LUT[28][9] ) );
  dp_1 \LUT_reg[28][8]  ( .ip(n13922), .ck(clk), .q(\LUT[28][8] ) );
  dp_1 \LUT_reg[28][7]  ( .ip(n13921), .ck(clk), .q(\LUT[28][7] ) );
  dp_1 \LUT_reg[28][6]  ( .ip(n13920), .ck(clk), .q(\LUT[28][6] ) );
  dp_1 \LUT_reg[28][5]  ( .ip(n13919), .ck(clk), .q(\LUT[28][5] ) );
  dp_1 \LUT_reg[28][4]  ( .ip(n13918), .ck(clk), .q(\LUT[28][4] ) );
  dp_1 \LUT_reg[28][3]  ( .ip(n13917), .ck(clk), .q(\LUT[28][3] ) );
  dp_1 \LUT_reg[28][2]  ( .ip(n13916), .ck(clk), .q(\LUT[28][2] ) );
  dp_1 \LUT_reg[28][1]  ( .ip(n13915), .ck(clk), .q(\LUT[28][1] ) );
  dp_1 \LUT_reg[28][0]  ( .ip(n13914), .ck(clk), .q(\LUT[28][0] ) );
  dp_1 \LUT_reg[27][15]  ( .ip(n13913), .ck(clk), .q(\LUT[27][15] ) );
  dp_1 \LUT_reg[27][14]  ( .ip(n13912), .ck(clk), .q(\LUT[27][14] ) );
  dp_1 \LUT_reg[27][13]  ( .ip(n13911), .ck(clk), .q(\LUT[27][13] ) );
  dp_1 \LUT_reg[27][12]  ( .ip(n13910), .ck(clk), .q(\LUT[27][12] ) );
  dp_1 \LUT_reg[27][11]  ( .ip(n13909), .ck(clk), .q(\LUT[27][11] ) );
  dp_1 \LUT_reg[27][10]  ( .ip(n13908), .ck(clk), .q(\LUT[27][10] ) );
  dp_1 \LUT_reg[27][9]  ( .ip(n13907), .ck(clk), .q(\LUT[27][9] ) );
  dp_1 \LUT_reg[27][8]  ( .ip(n13906), .ck(clk), .q(\LUT[27][8] ) );
  dp_1 \LUT_reg[27][7]  ( .ip(n13905), .ck(clk), .q(\LUT[27][7] ) );
  dp_1 \LUT_reg[27][6]  ( .ip(n13904), .ck(clk), .q(\LUT[27][6] ) );
  dp_1 \LUT_reg[27][5]  ( .ip(n13903), .ck(clk), .q(\LUT[27][5] ) );
  dp_1 \LUT_reg[27][4]  ( .ip(n13902), .ck(clk), .q(\LUT[27][4] ) );
  dp_1 \LUT_reg[27][3]  ( .ip(n13901), .ck(clk), .q(\LUT[27][3] ) );
  dp_1 \LUT_reg[27][2]  ( .ip(n13900), .ck(clk), .q(\LUT[27][2] ) );
  dp_1 \LUT_reg[27][1]  ( .ip(n13899), .ck(clk), .q(\LUT[27][1] ) );
  dp_1 \LUT_reg[27][0]  ( .ip(n13898), .ck(clk), .q(\LUT[27][0] ) );
  dp_1 \LUT_reg[26][15]  ( .ip(n13897), .ck(clk), .q(\LUT[26][15] ) );
  dp_1 \LUT_reg[26][14]  ( .ip(n13896), .ck(clk), .q(\LUT[26][14] ) );
  dp_1 \LUT_reg[26][13]  ( .ip(n13895), .ck(clk), .q(\LUT[26][13] ) );
  dp_1 \LUT_reg[26][12]  ( .ip(n13894), .ck(clk), .q(\LUT[26][12] ) );
  dp_1 \LUT_reg[26][11]  ( .ip(n13893), .ck(clk), .q(\LUT[26][11] ) );
  dp_1 \LUT_reg[26][10]  ( .ip(n13892), .ck(clk), .q(\LUT[26][10] ) );
  dp_1 \LUT_reg[26][9]  ( .ip(n13891), .ck(clk), .q(\LUT[26][9] ) );
  dp_1 \LUT_reg[26][8]  ( .ip(n13890), .ck(clk), .q(\LUT[26][8] ) );
  dp_1 \LUT_reg[26][7]  ( .ip(n13889), .ck(clk), .q(\LUT[26][7] ) );
  dp_1 \LUT_reg[26][6]  ( .ip(n13888), .ck(clk), .q(\LUT[26][6] ) );
  dp_1 \LUT_reg[26][5]  ( .ip(n13887), .ck(clk), .q(\LUT[26][5] ) );
  dp_1 \LUT_reg[26][4]  ( .ip(n13886), .ck(clk), .q(\LUT[26][4] ) );
  dp_1 \LUT_reg[26][3]  ( .ip(n13885), .ck(clk), .q(\LUT[26][3] ) );
  dp_1 \LUT_reg[26][2]  ( .ip(n13884), .ck(clk), .q(\LUT[26][2] ) );
  dp_1 \LUT_reg[26][1]  ( .ip(n13883), .ck(clk), .q(\LUT[26][1] ) );
  dp_1 \LUT_reg[26][0]  ( .ip(n13882), .ck(clk), .q(\LUT[26][0] ) );
  dp_1 \LUT_reg[25][15]  ( .ip(n13881), .ck(clk), .q(\LUT[25][15] ) );
  dp_1 \LUT_reg[25][14]  ( .ip(n13880), .ck(clk), .q(\LUT[25][14] ) );
  dp_1 \LUT_reg[25][13]  ( .ip(n13879), .ck(clk), .q(\LUT[25][13] ) );
  dp_1 \LUT_reg[25][12]  ( .ip(n13878), .ck(clk), .q(\LUT[25][12] ) );
  dp_1 \LUT_reg[25][11]  ( .ip(n13877), .ck(clk), .q(\LUT[25][11] ) );
  dp_1 \LUT_reg[25][10]  ( .ip(n13876), .ck(clk), .q(\LUT[25][10] ) );
  dp_1 \LUT_reg[25][9]  ( .ip(n13875), .ck(clk), .q(\LUT[25][9] ) );
  dp_1 \LUT_reg[25][8]  ( .ip(n13874), .ck(clk), .q(\LUT[25][8] ) );
  dp_1 \LUT_reg[25][7]  ( .ip(n13873), .ck(clk), .q(\LUT[25][7] ) );
  dp_1 \LUT_reg[25][6]  ( .ip(n13872), .ck(clk), .q(\LUT[25][6] ) );
  dp_1 \LUT_reg[25][5]  ( .ip(n13871), .ck(clk), .q(\LUT[25][5] ) );
  dp_1 \LUT_reg[25][4]  ( .ip(n13870), .ck(clk), .q(\LUT[25][4] ) );
  dp_1 \LUT_reg[25][3]  ( .ip(n13869), .ck(clk), .q(\LUT[25][3] ) );
  dp_1 \LUT_reg[25][2]  ( .ip(n13868), .ck(clk), .q(\LUT[25][2] ) );
  dp_1 \LUT_reg[25][1]  ( .ip(n13867), .ck(clk), .q(\LUT[25][1] ) );
  dp_1 \LUT_reg[25][0]  ( .ip(n13866), .ck(clk), .q(\LUT[25][0] ) );
  dp_1 \LUT_reg[24][15]  ( .ip(n13865), .ck(clk), .q(\LUT[24][15] ) );
  dp_1 \LUT_reg[24][14]  ( .ip(n13864), .ck(clk), .q(\LUT[24][14] ) );
  dp_1 \LUT_reg[24][13]  ( .ip(n13863), .ck(clk), .q(\LUT[24][13] ) );
  dp_1 \LUT_reg[24][12]  ( .ip(n13862), .ck(clk), .q(\LUT[24][12] ) );
  dp_1 \LUT_reg[24][11]  ( .ip(n13861), .ck(clk), .q(\LUT[24][11] ) );
  dp_1 \LUT_reg[24][10]  ( .ip(n13860), .ck(clk), .q(\LUT[24][10] ) );
  dp_1 \LUT_reg[24][9]  ( .ip(n13859), .ck(clk), .q(\LUT[24][9] ) );
  dp_1 \LUT_reg[24][8]  ( .ip(n13858), .ck(clk), .q(\LUT[24][8] ) );
  dp_1 \LUT_reg[24][7]  ( .ip(n13857), .ck(clk), .q(\LUT[24][7] ) );
  dp_1 \LUT_reg[24][6]  ( .ip(n13856), .ck(clk), .q(\LUT[24][6] ) );
  dp_1 \LUT_reg[24][5]  ( .ip(n13855), .ck(clk), .q(\LUT[24][5] ) );
  dp_1 \LUT_reg[24][4]  ( .ip(n13854), .ck(clk), .q(\LUT[24][4] ) );
  dp_1 \LUT_reg[24][3]  ( .ip(n13853), .ck(clk), .q(\LUT[24][3] ) );
  dp_1 \LUT_reg[24][2]  ( .ip(n13852), .ck(clk), .q(\LUT[24][2] ) );
  dp_1 \LUT_reg[24][1]  ( .ip(n13851), .ck(clk), .q(\LUT[24][1] ) );
  dp_1 \LUT_reg[24][0]  ( .ip(n13850), .ck(clk), .q(\LUT[24][0] ) );
  dp_1 \LUT_reg[23][15]  ( .ip(n13849), .ck(clk), .q(\LUT[23][15] ) );
  dp_1 \LUT_reg[23][14]  ( .ip(n13848), .ck(clk), .q(\LUT[23][14] ) );
  dp_1 \LUT_reg[23][13]  ( .ip(n13847), .ck(clk), .q(\LUT[23][13] ) );
  dp_1 \LUT_reg[23][12]  ( .ip(n13846), .ck(clk), .q(\LUT[23][12] ) );
  dp_1 \LUT_reg[23][11]  ( .ip(n13845), .ck(clk), .q(\LUT[23][11] ) );
  dp_1 \LUT_reg[23][10]  ( .ip(n13844), .ck(clk), .q(\LUT[23][10] ) );
  dp_1 \LUT_reg[23][9]  ( .ip(n13843), .ck(clk), .q(\LUT[23][9] ) );
  dp_1 \LUT_reg[23][8]  ( .ip(n13842), .ck(clk), .q(\LUT[23][8] ) );
  dp_1 \LUT_reg[23][7]  ( .ip(n13841), .ck(clk), .q(\LUT[23][7] ) );
  dp_1 \LUT_reg[23][6]  ( .ip(n13840), .ck(clk), .q(\LUT[23][6] ) );
  dp_1 \LUT_reg[23][5]  ( .ip(n13839), .ck(clk), .q(\LUT[23][5] ) );
  dp_1 \LUT_reg[23][4]  ( .ip(n13838), .ck(clk), .q(\LUT[23][4] ) );
  dp_1 \LUT_reg[23][3]  ( .ip(n13837), .ck(clk), .q(\LUT[23][3] ) );
  dp_1 \LUT_reg[23][2]  ( .ip(n13836), .ck(clk), .q(\LUT[23][2] ) );
  dp_1 \LUT_reg[23][1]  ( .ip(n13835), .ck(clk), .q(\LUT[23][1] ) );
  dp_1 \LUT_reg[23][0]  ( .ip(n13834), .ck(clk), .q(\LUT[23][0] ) );
  dp_1 \LUT_reg[22][15]  ( .ip(n13833), .ck(clk), .q(\LUT[22][15] ) );
  dp_1 \LUT_reg[22][14]  ( .ip(n13832), .ck(clk), .q(\LUT[22][14] ) );
  dp_1 \LUT_reg[22][13]  ( .ip(n13831), .ck(clk), .q(\LUT[22][13] ) );
  dp_1 \LUT_reg[22][12]  ( .ip(n13830), .ck(clk), .q(\LUT[22][12] ) );
  dp_1 \LUT_reg[22][11]  ( .ip(n13829), .ck(clk), .q(\LUT[22][11] ) );
  dp_1 \LUT_reg[22][10]  ( .ip(n13828), .ck(clk), .q(\LUT[22][10] ) );
  dp_1 \LUT_reg[22][9]  ( .ip(n13827), .ck(clk), .q(\LUT[22][9] ) );
  dp_1 \LUT_reg[22][8]  ( .ip(n13826), .ck(clk), .q(\LUT[22][8] ) );
  dp_1 \LUT_reg[22][7]  ( .ip(n13825), .ck(clk), .q(\LUT[22][7] ) );
  dp_1 \LUT_reg[22][6]  ( .ip(n13824), .ck(clk), .q(\LUT[22][6] ) );
  dp_1 \LUT_reg[22][5]  ( .ip(n13823), .ck(clk), .q(\LUT[22][5] ) );
  dp_1 \LUT_reg[22][4]  ( .ip(n13822), .ck(clk), .q(\LUT[22][4] ) );
  dp_1 \LUT_reg[22][3]  ( .ip(n13821), .ck(clk), .q(\LUT[22][3] ) );
  dp_1 \LUT_reg[22][2]  ( .ip(n13820), .ck(clk), .q(\LUT[22][2] ) );
  dp_1 \LUT_reg[22][1]  ( .ip(n13819), .ck(clk), .q(\LUT[22][1] ) );
  dp_1 \LUT_reg[22][0]  ( .ip(n13818), .ck(clk), .q(\LUT[22][0] ) );
  dp_1 \LUT_reg[21][15]  ( .ip(n13817), .ck(clk), .q(\LUT[21][15] ) );
  dp_1 \LUT_reg[21][14]  ( .ip(n13816), .ck(clk), .q(\LUT[21][14] ) );
  dp_1 \LUT_reg[21][13]  ( .ip(n13815), .ck(clk), .q(\LUT[21][13] ) );
  dp_1 \LUT_reg[21][12]  ( .ip(n13814), .ck(clk), .q(\LUT[21][12] ) );
  dp_1 \LUT_reg[21][11]  ( .ip(n13813), .ck(clk), .q(\LUT[21][11] ) );
  dp_1 \LUT_reg[21][10]  ( .ip(n13812), .ck(clk), .q(\LUT[21][10] ) );
  dp_1 \LUT_reg[21][9]  ( .ip(n13811), .ck(clk), .q(\LUT[21][9] ) );
  dp_1 \LUT_reg[21][8]  ( .ip(n13810), .ck(clk), .q(\LUT[21][8] ) );
  dp_1 \LUT_reg[21][7]  ( .ip(n13809), .ck(clk), .q(\LUT[21][7] ) );
  dp_1 \LUT_reg[21][6]  ( .ip(n13808), .ck(clk), .q(\LUT[21][6] ) );
  dp_1 \LUT_reg[21][5]  ( .ip(n13807), .ck(clk), .q(\LUT[21][5] ) );
  dp_1 \LUT_reg[21][4]  ( .ip(n13806), .ck(clk), .q(\LUT[21][4] ) );
  dp_1 \LUT_reg[21][3]  ( .ip(n13805), .ck(clk), .q(\LUT[21][3] ) );
  dp_1 \LUT_reg[21][2]  ( .ip(n13804), .ck(clk), .q(\LUT[21][2] ) );
  dp_1 \LUT_reg[21][1]  ( .ip(n13803), .ck(clk), .q(\LUT[21][1] ) );
  dp_1 \LUT_reg[21][0]  ( .ip(n13802), .ck(clk), .q(\LUT[21][0] ) );
  dp_1 \LUT_reg[20][15]  ( .ip(n13801), .ck(clk), .q(\LUT[20][15] ) );
  dp_1 \LUT_reg[20][14]  ( .ip(n13800), .ck(clk), .q(\LUT[20][14] ) );
  dp_1 \LUT_reg[20][13]  ( .ip(n13799), .ck(clk), .q(\LUT[20][13] ) );
  dp_1 \LUT_reg[20][12]  ( .ip(n13798), .ck(clk), .q(\LUT[20][12] ) );
  dp_1 \LUT_reg[20][11]  ( .ip(n13797), .ck(clk), .q(\LUT[20][11] ) );
  dp_1 \LUT_reg[20][10]  ( .ip(n13796), .ck(clk), .q(\LUT[20][10] ) );
  dp_1 \LUT_reg[20][9]  ( .ip(n13795), .ck(clk), .q(\LUT[20][9] ) );
  dp_1 \LUT_reg[20][8]  ( .ip(n13794), .ck(clk), .q(\LUT[20][8] ) );
  dp_1 \LUT_reg[20][7]  ( .ip(n13793), .ck(clk), .q(\LUT[20][7] ) );
  dp_1 \LUT_reg[20][6]  ( .ip(n13792), .ck(clk), .q(\LUT[20][6] ) );
  dp_1 \LUT_reg[20][5]  ( .ip(n13791), .ck(clk), .q(\LUT[20][5] ) );
  dp_1 \LUT_reg[20][4]  ( .ip(n13790), .ck(clk), .q(\LUT[20][4] ) );
  dp_1 \LUT_reg[20][3]  ( .ip(n13789), .ck(clk), .q(\LUT[20][3] ) );
  dp_1 \LUT_reg[20][2]  ( .ip(n13788), .ck(clk), .q(\LUT[20][2] ) );
  dp_1 \LUT_reg[20][1]  ( .ip(n13787), .ck(clk), .q(\LUT[20][1] ) );
  dp_1 \LUT_reg[20][0]  ( .ip(n13786), .ck(clk), .q(\LUT[20][0] ) );
  dp_1 \LUT_reg[19][15]  ( .ip(n13785), .ck(clk), .q(\LUT[19][15] ) );
  dp_1 \LUT_reg[19][14]  ( .ip(n13784), .ck(clk), .q(\LUT[19][14] ) );
  dp_1 \LUT_reg[19][13]  ( .ip(n13783), .ck(clk), .q(\LUT[19][13] ) );
  dp_1 \LUT_reg[19][12]  ( .ip(n13782), .ck(clk), .q(\LUT[19][12] ) );
  dp_1 \LUT_reg[19][11]  ( .ip(n13781), .ck(clk), .q(\LUT[19][11] ) );
  dp_1 \LUT_reg[19][10]  ( .ip(n13780), .ck(clk), .q(\LUT[19][10] ) );
  dp_1 \LUT_reg[19][9]  ( .ip(n13779), .ck(clk), .q(\LUT[19][9] ) );
  dp_1 \LUT_reg[19][8]  ( .ip(n13778), .ck(clk), .q(\LUT[19][8] ) );
  dp_1 \LUT_reg[19][7]  ( .ip(n13777), .ck(clk), .q(\LUT[19][7] ) );
  dp_1 \LUT_reg[19][6]  ( .ip(n13776), .ck(clk), .q(\LUT[19][6] ) );
  dp_1 \LUT_reg[19][5]  ( .ip(n13775), .ck(clk), .q(\LUT[19][5] ) );
  dp_1 \LUT_reg[19][4]  ( .ip(n13774), .ck(clk), .q(\LUT[19][4] ) );
  dp_1 \LUT_reg[19][3]  ( .ip(n13773), .ck(clk), .q(\LUT[19][3] ) );
  dp_1 \LUT_reg[19][2]  ( .ip(n13772), .ck(clk), .q(\LUT[19][2] ) );
  dp_1 \LUT_reg[19][1]  ( .ip(n13771), .ck(clk), .q(\LUT[19][1] ) );
  dp_1 \LUT_reg[19][0]  ( .ip(n13770), .ck(clk), .q(\LUT[19][0] ) );
  dp_1 \LUT_reg[18][15]  ( .ip(n13769), .ck(clk), .q(\LUT[18][15] ) );
  dp_1 \LUT_reg[18][14]  ( .ip(n13768), .ck(clk), .q(\LUT[18][14] ) );
  dp_1 \LUT_reg[18][13]  ( .ip(n13767), .ck(clk), .q(\LUT[18][13] ) );
  dp_1 \LUT_reg[18][12]  ( .ip(n13766), .ck(clk), .q(\LUT[18][12] ) );
  dp_1 \LUT_reg[18][11]  ( .ip(n13765), .ck(clk), .q(\LUT[18][11] ) );
  dp_1 \LUT_reg[18][10]  ( .ip(n13764), .ck(clk), .q(\LUT[18][10] ) );
  dp_1 \LUT_reg[18][9]  ( .ip(n13763), .ck(clk), .q(\LUT[18][9] ) );
  dp_1 \LUT_reg[18][8]  ( .ip(n13762), .ck(clk), .q(\LUT[18][8] ) );
  dp_1 \LUT_reg[18][7]  ( .ip(n13761), .ck(clk), .q(\LUT[18][7] ) );
  dp_1 \LUT_reg[18][6]  ( .ip(n13760), .ck(clk), .q(\LUT[18][6] ) );
  dp_1 \LUT_reg[18][5]  ( .ip(n13759), .ck(clk), .q(\LUT[18][5] ) );
  dp_1 \LUT_reg[18][4]  ( .ip(n13758), .ck(clk), .q(\LUT[18][4] ) );
  dp_1 \LUT_reg[18][3]  ( .ip(n13757), .ck(clk), .q(\LUT[18][3] ) );
  dp_1 \LUT_reg[18][2]  ( .ip(n13756), .ck(clk), .q(\LUT[18][2] ) );
  dp_1 \LUT_reg[18][1]  ( .ip(n13755), .ck(clk), .q(\LUT[18][1] ) );
  dp_1 \LUT_reg[18][0]  ( .ip(n13754), .ck(clk), .q(\LUT[18][0] ) );
  dp_1 \LUT_reg[17][15]  ( .ip(n13753), .ck(clk), .q(\LUT[17][15] ) );
  dp_1 \LUT_reg[17][14]  ( .ip(n13752), .ck(clk), .q(\LUT[17][14] ) );
  dp_1 \LUT_reg[17][13]  ( .ip(n13751), .ck(clk), .q(\LUT[17][13] ) );
  dp_1 \LUT_reg[17][12]  ( .ip(n13750), .ck(clk), .q(\LUT[17][12] ) );
  dp_1 \LUT_reg[17][11]  ( .ip(n13749), .ck(clk), .q(\LUT[17][11] ) );
  dp_1 \LUT_reg[17][10]  ( .ip(n13748), .ck(clk), .q(\LUT[17][10] ) );
  dp_1 \LUT_reg[17][9]  ( .ip(n13747), .ck(clk), .q(\LUT[17][9] ) );
  dp_1 \LUT_reg[17][8]  ( .ip(n13746), .ck(clk), .q(\LUT[17][8] ) );
  dp_1 \LUT_reg[17][7]  ( .ip(n13745), .ck(clk), .q(\LUT[17][7] ) );
  dp_1 \LUT_reg[17][6]  ( .ip(n13744), .ck(clk), .q(\LUT[17][6] ) );
  dp_1 \LUT_reg[17][5]  ( .ip(n13743), .ck(clk), .q(\LUT[17][5] ) );
  dp_1 \LUT_reg[17][4]  ( .ip(n13742), .ck(clk), .q(\LUT[17][4] ) );
  dp_1 \LUT_reg[17][3]  ( .ip(n13741), .ck(clk), .q(\LUT[17][3] ) );
  dp_1 \LUT_reg[17][2]  ( .ip(n13740), .ck(clk), .q(\LUT[17][2] ) );
  dp_1 \LUT_reg[17][1]  ( .ip(n13739), .ck(clk), .q(\LUT[17][1] ) );
  dp_1 \LUT_reg[17][0]  ( .ip(n13738), .ck(clk), .q(\LUT[17][0] ) );
  dp_1 \LUT_reg[16][15]  ( .ip(n13737), .ck(clk), .q(\LUT[16][15] ) );
  dp_1 \LUT_reg[16][14]  ( .ip(n13736), .ck(clk), .q(\LUT[16][14] ) );
  dp_1 \LUT_reg[16][13]  ( .ip(n13735), .ck(clk), .q(\LUT[16][13] ) );
  dp_1 \LUT_reg[16][12]  ( .ip(n13734), .ck(clk), .q(\LUT[16][12] ) );
  dp_1 \LUT_reg[16][11]  ( .ip(n13733), .ck(clk), .q(\LUT[16][11] ) );
  dp_1 \LUT_reg[16][10]  ( .ip(n13732), .ck(clk), .q(\LUT[16][10] ) );
  dp_1 \LUT_reg[16][9]  ( .ip(n13731), .ck(clk), .q(\LUT[16][9] ) );
  dp_1 \LUT_reg[16][8]  ( .ip(n13730), .ck(clk), .q(\LUT[16][8] ) );
  dp_1 \LUT_reg[16][7]  ( .ip(n13729), .ck(clk), .q(\LUT[16][7] ) );
  dp_1 \LUT_reg[16][6]  ( .ip(n13728), .ck(clk), .q(\LUT[16][6] ) );
  dp_1 \LUT_reg[16][5]  ( .ip(n13727), .ck(clk), .q(\LUT[16][5] ) );
  dp_1 \LUT_reg[16][4]  ( .ip(n13726), .ck(clk), .q(\LUT[16][4] ) );
  dp_1 \LUT_reg[16][3]  ( .ip(n13725), .ck(clk), .q(\LUT[16][3] ) );
  dp_1 \LUT_reg[16][2]  ( .ip(n13724), .ck(clk), .q(\LUT[16][2] ) );
  dp_1 \LUT_reg[16][1]  ( .ip(n13723), .ck(clk), .q(\LUT[16][1] ) );
  dp_1 \LUT_reg[16][0]  ( .ip(n13722), .ck(clk), .q(\LUT[16][0] ) );
  dp_1 \LUT_reg[15][15]  ( .ip(n13721), .ck(clk), .q(\LUT[15][15] ) );
  dp_1 \LUT_reg[15][14]  ( .ip(n13720), .ck(clk), .q(\LUT[15][14] ) );
  dp_1 \LUT_reg[15][13]  ( .ip(n13719), .ck(clk), .q(\LUT[15][13] ) );
  dp_1 \LUT_reg[15][12]  ( .ip(n13718), .ck(clk), .q(\LUT[15][12] ) );
  dp_1 \LUT_reg[15][11]  ( .ip(n13717), .ck(clk), .q(\LUT[15][11] ) );
  dp_1 \LUT_reg[15][10]  ( .ip(n13716), .ck(clk), .q(\LUT[15][10] ) );
  dp_1 \LUT_reg[15][9]  ( .ip(n13715), .ck(clk), .q(\LUT[15][9] ) );
  dp_1 \LUT_reg[15][8]  ( .ip(n13714), .ck(clk), .q(\LUT[15][8] ) );
  dp_1 \LUT_reg[15][7]  ( .ip(n13713), .ck(clk), .q(\LUT[15][7] ) );
  dp_1 \LUT_reg[15][6]  ( .ip(n13712), .ck(clk), .q(\LUT[15][6] ) );
  dp_1 \LUT_reg[15][5]  ( .ip(n13711), .ck(clk), .q(\LUT[15][5] ) );
  dp_1 \LUT_reg[15][4]  ( .ip(n13710), .ck(clk), .q(\LUT[15][4] ) );
  dp_1 \LUT_reg[15][3]  ( .ip(n13709), .ck(clk), .q(\LUT[15][3] ) );
  dp_1 \LUT_reg[15][2]  ( .ip(n13708), .ck(clk), .q(\LUT[15][2] ) );
  dp_1 \LUT_reg[15][1]  ( .ip(n13707), .ck(clk), .q(\LUT[15][1] ) );
  dp_1 \LUT_reg[15][0]  ( .ip(n13706), .ck(clk), .q(\LUT[15][0] ) );
  dp_1 \LUT_reg[14][15]  ( .ip(n13705), .ck(clk), .q(\LUT[14][15] ) );
  dp_1 \LUT_reg[14][14]  ( .ip(n13704), .ck(clk), .q(\LUT[14][14] ) );
  dp_1 \LUT_reg[14][13]  ( .ip(n13703), .ck(clk), .q(\LUT[14][13] ) );
  dp_1 \LUT_reg[14][12]  ( .ip(n13702), .ck(clk), .q(\LUT[14][12] ) );
  dp_1 \LUT_reg[14][11]  ( .ip(n13701), .ck(clk), .q(\LUT[14][11] ) );
  dp_1 \LUT_reg[14][10]  ( .ip(n13700), .ck(clk), .q(\LUT[14][10] ) );
  dp_1 \LUT_reg[14][9]  ( .ip(n13699), .ck(clk), .q(\LUT[14][9] ) );
  dp_1 \LUT_reg[14][8]  ( .ip(n13698), .ck(clk), .q(\LUT[14][8] ) );
  dp_1 \LUT_reg[14][7]  ( .ip(n13697), .ck(clk), .q(\LUT[14][7] ) );
  dp_1 \LUT_reg[14][6]  ( .ip(n13696), .ck(clk), .q(\LUT[14][6] ) );
  dp_1 \LUT_reg[14][5]  ( .ip(n13695), .ck(clk), .q(\LUT[14][5] ) );
  dp_1 \LUT_reg[14][4]  ( .ip(n13694), .ck(clk), .q(\LUT[14][4] ) );
  dp_1 \LUT_reg[14][3]  ( .ip(n13693), .ck(clk), .q(\LUT[14][3] ) );
  dp_1 \LUT_reg[14][2]  ( .ip(n13692), .ck(clk), .q(\LUT[14][2] ) );
  dp_1 \LUT_reg[14][1]  ( .ip(n13691), .ck(clk), .q(\LUT[14][1] ) );
  dp_1 \LUT_reg[14][0]  ( .ip(n13690), .ck(clk), .q(\LUT[14][0] ) );
  dp_1 \LUT_reg[13][15]  ( .ip(n13689), .ck(clk), .q(\LUT[13][15] ) );
  dp_1 \LUT_reg[13][14]  ( .ip(n13688), .ck(clk), .q(\LUT[13][14] ) );
  dp_1 \LUT_reg[13][13]  ( .ip(n13687), .ck(clk), .q(\LUT[13][13] ) );
  dp_1 \LUT_reg[13][12]  ( .ip(n13686), .ck(clk), .q(\LUT[13][12] ) );
  dp_1 \LUT_reg[13][11]  ( .ip(n13685), .ck(clk), .q(\LUT[13][11] ) );
  dp_1 \LUT_reg[13][10]  ( .ip(n13684), .ck(clk), .q(\LUT[13][10] ) );
  dp_1 \LUT_reg[13][9]  ( .ip(n13683), .ck(clk), .q(\LUT[13][9] ) );
  dp_1 \LUT_reg[13][8]  ( .ip(n13682), .ck(clk), .q(\LUT[13][8] ) );
  dp_1 \LUT_reg[13][7]  ( .ip(n13681), .ck(clk), .q(\LUT[13][7] ) );
  dp_1 \LUT_reg[13][6]  ( .ip(n13680), .ck(clk), .q(\LUT[13][6] ) );
  dp_1 \LUT_reg[13][5]  ( .ip(n13679), .ck(clk), .q(\LUT[13][5] ) );
  dp_1 \LUT_reg[13][4]  ( .ip(n13678), .ck(clk), .q(\LUT[13][4] ) );
  dp_1 \LUT_reg[13][3]  ( .ip(n13677), .ck(clk), .q(\LUT[13][3] ) );
  dp_1 \LUT_reg[13][2]  ( .ip(n13676), .ck(clk), .q(\LUT[13][2] ) );
  dp_1 \LUT_reg[13][1]  ( .ip(n13675), .ck(clk), .q(\LUT[13][1] ) );
  dp_1 \LUT_reg[13][0]  ( .ip(n13674), .ck(clk), .q(\LUT[13][0] ) );
  dp_1 \LUT_reg[12][15]  ( .ip(n13673), .ck(clk), .q(\LUT[12][15] ) );
  dp_1 \LUT_reg[12][14]  ( .ip(n13672), .ck(clk), .q(\LUT[12][14] ) );
  dp_1 \LUT_reg[12][13]  ( .ip(n13671), .ck(clk), .q(\LUT[12][13] ) );
  dp_1 \LUT_reg[12][12]  ( .ip(n13670), .ck(clk), .q(\LUT[12][12] ) );
  dp_1 \LUT_reg[12][11]  ( .ip(n13669), .ck(clk), .q(\LUT[12][11] ) );
  dp_1 \LUT_reg[12][10]  ( .ip(n13668), .ck(clk), .q(\LUT[12][10] ) );
  dp_1 \LUT_reg[12][9]  ( .ip(n13667), .ck(clk), .q(\LUT[12][9] ) );
  dp_1 \LUT_reg[12][8]  ( .ip(n13666), .ck(clk), .q(\LUT[12][8] ) );
  dp_1 \LUT_reg[12][7]  ( .ip(n13665), .ck(clk), .q(\LUT[12][7] ) );
  dp_1 \LUT_reg[12][6]  ( .ip(n13664), .ck(clk), .q(\LUT[12][6] ) );
  dp_1 \LUT_reg[12][5]  ( .ip(n13663), .ck(clk), .q(\LUT[12][5] ) );
  dp_1 \LUT_reg[12][4]  ( .ip(n13662), .ck(clk), .q(\LUT[12][4] ) );
  dp_1 \LUT_reg[12][3]  ( .ip(n13661), .ck(clk), .q(\LUT[12][3] ) );
  dp_1 \LUT_reg[12][2]  ( .ip(n13660), .ck(clk), .q(\LUT[12][2] ) );
  dp_1 \LUT_reg[12][1]  ( .ip(n13659), .ck(clk), .q(\LUT[12][1] ) );
  dp_1 \LUT_reg[12][0]  ( .ip(n13658), .ck(clk), .q(\LUT[12][0] ) );
  dp_1 \LUT_reg[11][15]  ( .ip(n13657), .ck(clk), .q(\LUT[11][15] ) );
  dp_1 \LUT_reg[11][14]  ( .ip(n13656), .ck(clk), .q(\LUT[11][14] ) );
  dp_1 \LUT_reg[11][13]  ( .ip(n13655), .ck(clk), .q(\LUT[11][13] ) );
  dp_1 \LUT_reg[11][12]  ( .ip(n13654), .ck(clk), .q(\LUT[11][12] ) );
  dp_1 \LUT_reg[11][11]  ( .ip(n13653), .ck(clk), .q(\LUT[11][11] ) );
  dp_1 \LUT_reg[11][10]  ( .ip(n13652), .ck(clk), .q(\LUT[11][10] ) );
  dp_1 \LUT_reg[11][9]  ( .ip(n13651), .ck(clk), .q(\LUT[11][9] ) );
  dp_1 \LUT_reg[11][8]  ( .ip(n13650), .ck(clk), .q(\LUT[11][8] ) );
  dp_1 \LUT_reg[11][7]  ( .ip(n13649), .ck(clk), .q(\LUT[11][7] ) );
  dp_1 \LUT_reg[11][6]  ( .ip(n13648), .ck(clk), .q(\LUT[11][6] ) );
  dp_1 \LUT_reg[11][5]  ( .ip(n13647), .ck(clk), .q(\LUT[11][5] ) );
  dp_1 \LUT_reg[11][4]  ( .ip(n13646), .ck(clk), .q(\LUT[11][4] ) );
  dp_1 \LUT_reg[11][3]  ( .ip(n13645), .ck(clk), .q(\LUT[11][3] ) );
  dp_1 \LUT_reg[11][2]  ( .ip(n13644), .ck(clk), .q(\LUT[11][2] ) );
  dp_1 \LUT_reg[11][1]  ( .ip(n13643), .ck(clk), .q(\LUT[11][1] ) );
  dp_1 \LUT_reg[11][0]  ( .ip(n13642), .ck(clk), .q(\LUT[11][0] ) );
  dp_1 \LUT_reg[10][15]  ( .ip(n13641), .ck(clk), .q(\LUT[10][15] ) );
  dp_1 \LUT_reg[10][14]  ( .ip(n13640), .ck(clk), .q(\LUT[10][14] ) );
  dp_1 \LUT_reg[10][13]  ( .ip(n13639), .ck(clk), .q(\LUT[10][13] ) );
  dp_1 \LUT_reg[10][12]  ( .ip(n13638), .ck(clk), .q(\LUT[10][12] ) );
  dp_1 \LUT_reg[10][11]  ( .ip(n13637), .ck(clk), .q(\LUT[10][11] ) );
  dp_1 \LUT_reg[10][10]  ( .ip(n13636), .ck(clk), .q(\LUT[10][10] ) );
  dp_1 \LUT_reg[10][9]  ( .ip(n13635), .ck(clk), .q(\LUT[10][9] ) );
  dp_1 \LUT_reg[10][8]  ( .ip(n13634), .ck(clk), .q(\LUT[10][8] ) );
  dp_1 \LUT_reg[10][7]  ( .ip(n13633), .ck(clk), .q(\LUT[10][7] ) );
  dp_1 \LUT_reg[10][6]  ( .ip(n13632), .ck(clk), .q(\LUT[10][6] ) );
  dp_1 \LUT_reg[10][5]  ( .ip(n13631), .ck(clk), .q(\LUT[10][5] ) );
  dp_1 \LUT_reg[10][4]  ( .ip(n13630), .ck(clk), .q(\LUT[10][4] ) );
  dp_1 \LUT_reg[10][3]  ( .ip(n13629), .ck(clk), .q(\LUT[10][3] ) );
  dp_1 \LUT_reg[10][2]  ( .ip(n13628), .ck(clk), .q(\LUT[10][2] ) );
  dp_1 \LUT_reg[10][1]  ( .ip(n13627), .ck(clk), .q(\LUT[10][1] ) );
  dp_1 \LUT_reg[10][0]  ( .ip(n13626), .ck(clk), .q(\LUT[10][0] ) );
  dp_1 \LUT_reg[9][15]  ( .ip(n13625), .ck(clk), .q(\LUT[9][15] ) );
  dp_1 \LUT_reg[9][14]  ( .ip(n13624), .ck(clk), .q(\LUT[9][14] ) );
  dp_1 \LUT_reg[9][13]  ( .ip(n13623), .ck(clk), .q(\LUT[9][13] ) );
  dp_1 \LUT_reg[9][12]  ( .ip(n13622), .ck(clk), .q(\LUT[9][12] ) );
  dp_1 \LUT_reg[9][11]  ( .ip(n13621), .ck(clk), .q(\LUT[9][11] ) );
  dp_1 \LUT_reg[9][10]  ( .ip(n13620), .ck(clk), .q(\LUT[9][10] ) );
  dp_1 \LUT_reg[9][9]  ( .ip(n13619), .ck(clk), .q(\LUT[9][9] ) );
  dp_1 \LUT_reg[9][8]  ( .ip(n13618), .ck(clk), .q(\LUT[9][8] ) );
  dp_1 \LUT_reg[9][7]  ( .ip(n13617), .ck(clk), .q(\LUT[9][7] ) );
  dp_1 \LUT_reg[9][6]  ( .ip(n13616), .ck(clk), .q(\LUT[9][6] ) );
  dp_1 \LUT_reg[9][5]  ( .ip(n13615), .ck(clk), .q(\LUT[9][5] ) );
  dp_1 \LUT_reg[9][4]  ( .ip(n13614), .ck(clk), .q(\LUT[9][4] ) );
  dp_1 \LUT_reg[9][3]  ( .ip(n13613), .ck(clk), .q(\LUT[9][3] ) );
  dp_1 \LUT_reg[9][2]  ( .ip(n13612), .ck(clk), .q(\LUT[9][2] ) );
  dp_1 \LUT_reg[9][1]  ( .ip(n13611), .ck(clk), .q(\LUT[9][1] ) );
  dp_1 \LUT_reg[9][0]  ( .ip(n13610), .ck(clk), .q(\LUT[9][0] ) );
  dp_1 \LUT_reg[8][15]  ( .ip(n13609), .ck(clk), .q(\LUT[8][15] ) );
  dp_1 \LUT_reg[8][14]  ( .ip(n13608), .ck(clk), .q(\LUT[8][14] ) );
  dp_1 \LUT_reg[8][13]  ( .ip(n13607), .ck(clk), .q(\LUT[8][13] ) );
  dp_1 \LUT_reg[8][12]  ( .ip(n13606), .ck(clk), .q(\LUT[8][12] ) );
  dp_1 \LUT_reg[8][11]  ( .ip(n13605), .ck(clk), .q(\LUT[8][11] ) );
  dp_1 \LUT_reg[8][10]  ( .ip(n13604), .ck(clk), .q(\LUT[8][10] ) );
  dp_1 \LUT_reg[8][9]  ( .ip(n13603), .ck(clk), .q(\LUT[8][9] ) );
  dp_1 \LUT_reg[8][8]  ( .ip(n13602), .ck(clk), .q(\LUT[8][8] ) );
  dp_1 \LUT_reg[8][7]  ( .ip(n13601), .ck(clk), .q(\LUT[8][7] ) );
  dp_1 \LUT_reg[8][6]  ( .ip(n13600), .ck(clk), .q(\LUT[8][6] ) );
  dp_1 \LUT_reg[8][5]  ( .ip(n13599), .ck(clk), .q(\LUT[8][5] ) );
  dp_1 \LUT_reg[8][4]  ( .ip(n13598), .ck(clk), .q(\LUT[8][4] ) );
  dp_1 \LUT_reg[8][3]  ( .ip(n13597), .ck(clk), .q(\LUT[8][3] ) );
  dp_1 \LUT_reg[8][2]  ( .ip(n13596), .ck(clk), .q(\LUT[8][2] ) );
  dp_1 \LUT_reg[8][1]  ( .ip(n13595), .ck(clk), .q(\LUT[8][1] ) );
  dp_1 \LUT_reg[8][0]  ( .ip(n13594), .ck(clk), .q(\LUT[8][0] ) );
  dp_1 \LUT_reg[7][15]  ( .ip(n13593), .ck(clk), .q(\LUT[7][15] ) );
  dp_1 \LUT_reg[7][14]  ( .ip(n13592), .ck(clk), .q(\LUT[7][14] ) );
  dp_1 \LUT_reg[7][13]  ( .ip(n13591), .ck(clk), .q(\LUT[7][13] ) );
  dp_1 \LUT_reg[7][12]  ( .ip(n13590), .ck(clk), .q(\LUT[7][12] ) );
  dp_1 \LUT_reg[7][11]  ( .ip(n13589), .ck(clk), .q(\LUT[7][11] ) );
  dp_1 \LUT_reg[7][10]  ( .ip(n13588), .ck(clk), .q(\LUT[7][10] ) );
  dp_1 \LUT_reg[7][9]  ( .ip(n13587), .ck(clk), .q(\LUT[7][9] ) );
  dp_1 \LUT_reg[7][8]  ( .ip(n13586), .ck(clk), .q(\LUT[7][8] ) );
  dp_1 \LUT_reg[7][7]  ( .ip(n13585), .ck(clk), .q(\LUT[7][7] ) );
  dp_1 \LUT_reg[7][6]  ( .ip(n13584), .ck(clk), .q(\LUT[7][6] ) );
  dp_1 \LUT_reg[7][5]  ( .ip(n13583), .ck(clk), .q(\LUT[7][5] ) );
  dp_1 \LUT_reg[7][4]  ( .ip(n13582), .ck(clk), .q(\LUT[7][4] ) );
  dp_1 \LUT_reg[7][3]  ( .ip(n13581), .ck(clk), .q(\LUT[7][3] ) );
  dp_1 \LUT_reg[7][2]  ( .ip(n13580), .ck(clk), .q(\LUT[7][2] ) );
  dp_1 \LUT_reg[7][1]  ( .ip(n13579), .ck(clk), .q(\LUT[7][1] ) );
  dp_1 \LUT_reg[7][0]  ( .ip(n13578), .ck(clk), .q(\LUT[7][0] ) );
  dp_1 \LUT_reg[6][15]  ( .ip(n13577), .ck(clk), .q(\LUT[6][15] ) );
  dp_1 \LUT_reg[6][14]  ( .ip(n13576), .ck(clk), .q(\LUT[6][14] ) );
  dp_1 \LUT_reg[6][13]  ( .ip(n13575), .ck(clk), .q(\LUT[6][13] ) );
  dp_1 \LUT_reg[6][12]  ( .ip(n13574), .ck(clk), .q(\LUT[6][12] ) );
  dp_1 \LUT_reg[6][11]  ( .ip(n13573), .ck(clk), .q(\LUT[6][11] ) );
  dp_1 \LUT_reg[6][10]  ( .ip(n13572), .ck(clk), .q(\LUT[6][10] ) );
  dp_1 \LUT_reg[6][9]  ( .ip(n13571), .ck(clk), .q(\LUT[6][9] ) );
  dp_1 \LUT_reg[6][8]  ( .ip(n13570), .ck(clk), .q(\LUT[6][8] ) );
  dp_1 \LUT_reg[6][7]  ( .ip(n13569), .ck(clk), .q(\LUT[6][7] ) );
  dp_1 \LUT_reg[6][6]  ( .ip(n13568), .ck(clk), .q(\LUT[6][6] ) );
  dp_1 \LUT_reg[6][5]  ( .ip(n13567), .ck(clk), .q(\LUT[6][5] ) );
  dp_1 \LUT_reg[6][4]  ( .ip(n13566), .ck(clk), .q(\LUT[6][4] ) );
  dp_1 \LUT_reg[6][3]  ( .ip(n13565), .ck(clk), .q(\LUT[6][3] ) );
  dp_1 \LUT_reg[6][2]  ( .ip(n13564), .ck(clk), .q(\LUT[6][2] ) );
  dp_1 \LUT_reg[6][1]  ( .ip(n13563), .ck(clk), .q(\LUT[6][1] ) );
  dp_1 \LUT_reg[6][0]  ( .ip(n13562), .ck(clk), .q(\LUT[6][0] ) );
  dp_1 \LUT_reg[5][15]  ( .ip(n13561), .ck(clk), .q(\LUT[5][15] ) );
  dp_1 \LUT_reg[5][14]  ( .ip(n13560), .ck(clk), .q(\LUT[5][14] ) );
  dp_1 \LUT_reg[5][13]  ( .ip(n13559), .ck(clk), .q(\LUT[5][13] ) );
  dp_1 \LUT_reg[5][12]  ( .ip(n13558), .ck(clk), .q(\LUT[5][12] ) );
  dp_1 \LUT_reg[5][11]  ( .ip(n13557), .ck(clk), .q(\LUT[5][11] ) );
  dp_1 \LUT_reg[5][10]  ( .ip(n13556), .ck(clk), .q(\LUT[5][10] ) );
  dp_1 \LUT_reg[5][9]  ( .ip(n13555), .ck(clk), .q(\LUT[5][9] ) );
  dp_1 \LUT_reg[5][8]  ( .ip(n13554), .ck(clk), .q(\LUT[5][8] ) );
  dp_1 \LUT_reg[5][7]  ( .ip(n13553), .ck(clk), .q(\LUT[5][7] ) );
  dp_1 \LUT_reg[5][6]  ( .ip(n13552), .ck(clk), .q(\LUT[5][6] ) );
  dp_1 \LUT_reg[5][5]  ( .ip(n13551), .ck(clk), .q(\LUT[5][5] ) );
  dp_1 \LUT_reg[5][4]  ( .ip(n13550), .ck(clk), .q(\LUT[5][4] ) );
  dp_1 \LUT_reg[5][3]  ( .ip(n13549), .ck(clk), .q(\LUT[5][3] ) );
  dp_1 \LUT_reg[5][2]  ( .ip(n13548), .ck(clk), .q(\LUT[5][2] ) );
  dp_1 \LUT_reg[5][1]  ( .ip(n13547), .ck(clk), .q(\LUT[5][1] ) );
  dp_1 \LUT_reg[5][0]  ( .ip(n13546), .ck(clk), .q(\LUT[5][0] ) );
  dp_1 \LUT_reg[4][15]  ( .ip(n13545), .ck(clk), .q(\LUT[4][15] ) );
  dp_1 \LUT_reg[4][14]  ( .ip(n13544), .ck(clk), .q(\LUT[4][14] ) );
  dp_1 \LUT_reg[4][13]  ( .ip(n13543), .ck(clk), .q(\LUT[4][13] ) );
  dp_1 \LUT_reg[4][12]  ( .ip(n13542), .ck(clk), .q(\LUT[4][12] ) );
  dp_1 \LUT_reg[4][11]  ( .ip(n13541), .ck(clk), .q(\LUT[4][11] ) );
  dp_1 \LUT_reg[4][10]  ( .ip(n13540), .ck(clk), .q(\LUT[4][10] ) );
  dp_1 \LUT_reg[4][9]  ( .ip(n13539), .ck(clk), .q(\LUT[4][9] ) );
  dp_1 \LUT_reg[4][8]  ( .ip(n13538), .ck(clk), .q(\LUT[4][8] ) );
  dp_1 \LUT_reg[4][7]  ( .ip(n13537), .ck(clk), .q(\LUT[4][7] ) );
  dp_1 \LUT_reg[4][6]  ( .ip(n13536), .ck(clk), .q(\LUT[4][6] ) );
  dp_1 \LUT_reg[4][5]  ( .ip(n13535), .ck(clk), .q(\LUT[4][5] ) );
  dp_1 \LUT_reg[4][4]  ( .ip(n13534), .ck(clk), .q(\LUT[4][4] ) );
  dp_1 \LUT_reg[4][3]  ( .ip(n13533), .ck(clk), .q(\LUT[4][3] ) );
  dp_1 \LUT_reg[4][2]  ( .ip(n13532), .ck(clk), .q(\LUT[4][2] ) );
  dp_1 \LUT_reg[4][1]  ( .ip(n13531), .ck(clk), .q(\LUT[4][1] ) );
  dp_1 \LUT_reg[4][0]  ( .ip(n13530), .ck(clk), .q(\LUT[4][0] ) );
  dp_1 \LUT_reg[3][15]  ( .ip(n13529), .ck(clk), .q(\LUT[3][15] ) );
  dp_1 \LUT_reg[3][14]  ( .ip(n13528), .ck(clk), .q(\LUT[3][14] ) );
  dp_1 \LUT_reg[3][13]  ( .ip(n13527), .ck(clk), .q(\LUT[3][13] ) );
  dp_1 \LUT_reg[3][12]  ( .ip(n13526), .ck(clk), .q(\LUT[3][12] ) );
  dp_1 \LUT_reg[3][11]  ( .ip(n13525), .ck(clk), .q(\LUT[3][11] ) );
  dp_1 \LUT_reg[3][10]  ( .ip(n13524), .ck(clk), .q(\LUT[3][10] ) );
  dp_1 \LUT_reg[3][9]  ( .ip(n13523), .ck(clk), .q(\LUT[3][9] ) );
  dp_1 \LUT_reg[3][8]  ( .ip(n13522), .ck(clk), .q(\LUT[3][8] ) );
  dp_1 \LUT_reg[3][7]  ( .ip(n13521), .ck(clk), .q(\LUT[3][7] ) );
  dp_1 \LUT_reg[3][6]  ( .ip(n13520), .ck(clk), .q(\LUT[3][6] ) );
  dp_1 \LUT_reg[3][5]  ( .ip(n13519), .ck(clk), .q(\LUT[3][5] ) );
  dp_1 \LUT_reg[3][4]  ( .ip(n13518), .ck(clk), .q(\LUT[3][4] ) );
  dp_1 \LUT_reg[3][3]  ( .ip(n13517), .ck(clk), .q(\LUT[3][3] ) );
  dp_1 \LUT_reg[3][2]  ( .ip(n13516), .ck(clk), .q(\LUT[3][2] ) );
  dp_1 \LUT_reg[3][1]  ( .ip(n13515), .ck(clk), .q(\LUT[3][1] ) );
  dp_1 \LUT_reg[3][0]  ( .ip(n13514), .ck(clk), .q(\LUT[3][0] ) );
  dp_1 \LUT_reg[2][15]  ( .ip(n13513), .ck(clk), .q(\LUT[2][15] ) );
  dp_1 \LUT_reg[2][14]  ( .ip(n13512), .ck(clk), .q(\LUT[2][14] ) );
  dp_1 \LUT_reg[2][13]  ( .ip(n13511), .ck(clk), .q(\LUT[2][13] ) );
  dp_1 \LUT_reg[2][12]  ( .ip(n13510), .ck(clk), .q(\LUT[2][12] ) );
  dp_1 \LUT_reg[2][11]  ( .ip(n13509), .ck(clk), .q(\LUT[2][11] ) );
  dp_1 \LUT_reg[2][10]  ( .ip(n13508), .ck(clk), .q(\LUT[2][10] ) );
  dp_1 \LUT_reg[2][9]  ( .ip(n13507), .ck(clk), .q(\LUT[2][9] ) );
  dp_1 \LUT_reg[2][8]  ( .ip(n13506), .ck(clk), .q(\LUT[2][8] ) );
  dp_1 \LUT_reg[2][7]  ( .ip(n13505), .ck(clk), .q(\LUT[2][7] ) );
  dp_1 \LUT_reg[2][6]  ( .ip(n13504), .ck(clk), .q(\LUT[2][6] ) );
  dp_1 \LUT_reg[2][5]  ( .ip(n13503), .ck(clk), .q(\LUT[2][5] ) );
  dp_1 \LUT_reg[2][4]  ( .ip(n13502), .ck(clk), .q(\LUT[2][4] ) );
  dp_1 \LUT_reg[2][3]  ( .ip(n13501), .ck(clk), .q(\LUT[2][3] ) );
  dp_1 \LUT_reg[2][2]  ( .ip(n13500), .ck(clk), .q(\LUT[2][2] ) );
  dp_1 \LUT_reg[2][1]  ( .ip(n13499), .ck(clk), .q(\LUT[2][1] ) );
  dp_1 \LUT_reg[2][0]  ( .ip(n13498), .ck(clk), .q(\LUT[2][0] ) );
  dp_1 \LUT_reg[1][15]  ( .ip(n13497), .ck(clk), .q(\LUT[1][15] ) );
  dp_1 \LUT_reg[1][14]  ( .ip(n13496), .ck(clk), .q(\LUT[1][14] ) );
  dp_1 \LUT_reg[1][13]  ( .ip(n13495), .ck(clk), .q(\LUT[1][13] ) );
  dp_1 \LUT_reg[1][12]  ( .ip(n13494), .ck(clk), .q(\LUT[1][12] ) );
  dp_1 \LUT_reg[1][11]  ( .ip(n13493), .ck(clk), .q(\LUT[1][11] ) );
  dp_1 \LUT_reg[1][10]  ( .ip(n13492), .ck(clk), .q(\LUT[1][10] ) );
  dp_1 \LUT_reg[1][9]  ( .ip(n13491), .ck(clk), .q(\LUT[1][9] ) );
  dp_1 \LUT_reg[1][8]  ( .ip(n13490), .ck(clk), .q(\LUT[1][8] ) );
  dp_1 \LUT_reg[1][7]  ( .ip(n13489), .ck(clk), .q(\LUT[1][7] ) );
  dp_1 \LUT_reg[1][6]  ( .ip(n13488), .ck(clk), .q(\LUT[1][6] ) );
  dp_1 \LUT_reg[1][5]  ( .ip(n13487), .ck(clk), .q(\LUT[1][5] ) );
  dp_1 \LUT_reg[1][4]  ( .ip(n13486), .ck(clk), .q(\LUT[1][4] ) );
  dp_1 \LUT_reg[1][3]  ( .ip(n13485), .ck(clk), .q(\LUT[1][3] ) );
  dp_1 \LUT_reg[1][2]  ( .ip(n13484), .ck(clk), .q(\LUT[1][2] ) );
  dp_1 \LUT_reg[1][1]  ( .ip(n13483), .ck(clk), .q(\LUT[1][1] ) );
  dp_1 \LUT_reg[1][0]  ( .ip(n13482), .ck(clk), .q(\LUT[1][0] ) );
  dp_1 \LUT_reg[0][15]  ( .ip(n13481), .ck(clk), .q(\LUT[0][15] ) );
  dp_1 \y_reg[15]  ( .ip(n13450), .ck(clk), .q(sig_out[15]) );
  dp_1 \LUT_reg[0][14]  ( .ip(n13480), .ck(clk), .q(\LUT[0][14] ) );
  dp_1 \y_reg[14]  ( .ip(n13451), .ck(clk), .q(sig_out[14]) );
  dp_1 \LUT_reg[0][13]  ( .ip(n13479), .ck(clk), .q(\LUT[0][13] ) );
  dp_1 \y_reg[13]  ( .ip(n13452), .ck(clk), .q(sig_out[13]) );
  dp_1 \LUT_reg[0][12]  ( .ip(n13478), .ck(clk), .q(\LUT[0][12] ) );
  dp_1 \y_reg[12]  ( .ip(n13453), .ck(clk), .q(sig_out[12]) );
  dp_1 \LUT_reg[0][11]  ( .ip(n13477), .ck(clk), .q(\LUT[0][11] ) );
  dp_1 \y_reg[11]  ( .ip(n13454), .ck(clk), .q(sig_out[11]) );
  dp_1 \LUT_reg[0][10]  ( .ip(n13476), .ck(clk), .q(\LUT[0][10] ) );
  dp_1 \y_reg[10]  ( .ip(n13455), .ck(clk), .q(sig_out[10]) );
  dp_1 \LUT_reg[0][9]  ( .ip(n13475), .ck(clk), .q(\LUT[0][9] ) );
  dp_1 \y_reg[9]  ( .ip(n13456), .ck(clk), .q(sig_out[9]) );
  dp_1 \LUT_reg[0][8]  ( .ip(n13474), .ck(clk), .q(\LUT[0][8] ) );
  dp_1 \y_reg[8]  ( .ip(n13457), .ck(clk), .q(sig_out[8]) );
  dp_1 \LUT_reg[0][7]  ( .ip(n13473), .ck(clk), .q(\LUT[0][7] ) );
  dp_1 \y_reg[7]  ( .ip(n13458), .ck(clk), .q(sig_out[7]) );
  dp_1 \LUT_reg[0][6]  ( .ip(n13472), .ck(clk), .q(\LUT[0][6] ) );
  dp_1 \y_reg[6]  ( .ip(n13459), .ck(clk), .q(sig_out[6]) );
  dp_1 \LUT_reg[0][5]  ( .ip(n13471), .ck(clk), .q(\LUT[0][5] ) );
  dp_1 \y_reg[5]  ( .ip(n13460), .ck(clk), .q(sig_out[5]) );
  dp_1 \LUT_reg[0][4]  ( .ip(n13470), .ck(clk), .q(\LUT[0][4] ) );
  dp_1 \y_reg[4]  ( .ip(n13461), .ck(clk), .q(sig_out[4]) );
  dp_1 \LUT_reg[0][3]  ( .ip(n13469), .ck(clk), .q(\LUT[0][3] ) );
  dp_1 \y_reg[3]  ( .ip(n13462), .ck(clk), .q(sig_out[3]) );
  dp_1 \LUT_reg[0][2]  ( .ip(n13468), .ck(clk), .q(\LUT[0][2] ) );
  dp_1 \y_reg[2]  ( .ip(n13463), .ck(clk), .q(sig_out[2]) );
  dp_1 \LUT_reg[0][1]  ( .ip(n13467), .ck(clk), .q(\LUT[0][1] ) );
  dp_1 \y_reg[1]  ( .ip(n13464), .ck(clk), .q(sig_out[1]) );
  dp_1 \LUT_reg[0][0]  ( .ip(n13466), .ck(clk), .q(\LUT[0][0] ) );
  dp_1 \y_reg[0]  ( .ip(n13465), .ck(clk), .q(sig_out[0]) );
  buf_1 U17324 ( .ip(d[15]), .op(n17333) );
  nor2_1 U17325 ( .ip1(address[2]), .ip2(address[1]), .op(n17331) );
  inv_1 U17326 ( .ip(address[3]), .op(n17324) );
  nor2_1 U17327 ( .ip1(address[0]), .ip2(n17324), .op(n17330) );
  nand2_1 U17328 ( .ip1(n17331), .ip2(n17330), .op(n17396) );
  nand4_1 U17329 ( .ip1(we), .ip2(address[4]), .ip3(address[6]), .ip4(
        address[5]), .op(n17326) );
  nor2_1 U17330 ( .ip1(n17396), .ip2(n17326), .op(n17323) );
  mux2_1 U17331 ( .ip1(\x[120][15] ), .ip2(n17333), .s(n17323), .op(n17322) );
  buf_1 U17332 ( .ip(d[14]), .op(n17334) );
  mux2_1 U17333 ( .ip1(\x[120][14] ), .ip2(n17334), .s(n17323), .op(n17321) );
  buf_1 U17334 ( .ip(d[13]), .op(n17335) );
  mux2_1 U17335 ( .ip1(\x[120][13] ), .ip2(n17335), .s(n17323), .op(n17320) );
  buf_1 U17336 ( .ip(d[12]), .op(n17336) );
  mux2_1 U17337 ( .ip1(\x[120][12] ), .ip2(n17336), .s(n17323), .op(n17319) );
  buf_1 U17338 ( .ip(d[11]), .op(n17337) );
  mux2_1 U17339 ( .ip1(\x[120][11] ), .ip2(n17337), .s(n17323), .op(n17318) );
  buf_1 U17340 ( .ip(d[10]), .op(n17338) );
  mux2_1 U17341 ( .ip1(\x[120][10] ), .ip2(n17338), .s(n17323), .op(n17317) );
  buf_1 U17342 ( .ip(d[9]), .op(n17339) );
  mux2_1 U17343 ( .ip1(\x[120][9] ), .ip2(n17339), .s(n17323), .op(n17316) );
  buf_1 U17344 ( .ip(d[8]), .op(n17340) );
  mux2_1 U17345 ( .ip1(\x[120][8] ), .ip2(n17340), .s(n17323), .op(n17315) );
  buf_1 U17346 ( .ip(d[7]), .op(n17341) );
  mux2_1 U17347 ( .ip1(\x[120][7] ), .ip2(n17341), .s(n17323), .op(n17314) );
  buf_1 U17348 ( .ip(d[6]), .op(n17342) );
  mux2_1 U17349 ( .ip1(\x[120][6] ), .ip2(n17342), .s(n17323), .op(n17313) );
  buf_1 U17350 ( .ip(d[5]), .op(n17343) );
  mux2_1 U17351 ( .ip1(\x[120][5] ), .ip2(n17343), .s(n17323), .op(n17312) );
  buf_1 U17352 ( .ip(d[4]), .op(n17344) );
  mux2_1 U17353 ( .ip1(\x[120][4] ), .ip2(n17344), .s(n17323), .op(n17311) );
  buf_1 U17354 ( .ip(d[3]), .op(n17345) );
  mux2_1 U17355 ( .ip1(\x[120][3] ), .ip2(n17345), .s(n17323), .op(n17310) );
  buf_1 U17356 ( .ip(d[2]), .op(n17346) );
  mux2_1 U17357 ( .ip1(\x[120][2] ), .ip2(n17346), .s(n17323), .op(n17309) );
  buf_1 U17358 ( .ip(d[1]), .op(n17347) );
  mux2_1 U17359 ( .ip1(\x[120][1] ), .ip2(n17347), .s(n17323), .op(n17308) );
  buf_1 U17360 ( .ip(d[0]), .op(n17348) );
  mux2_1 U17361 ( .ip1(\x[120][0] ), .ip2(n17348), .s(n17323), .op(n17307) );
  nand4_1 U17362 ( .ip1(address[1]), .ip2(address[2]), .ip3(address[0]), .ip4(
        n17324), .op(n17397) );
  nor2_1 U17363 ( .ip1(n17326), .ip2(n17397), .op(n17410) );
  mux2_1 U17364 ( .ip1(\x[119][15] ), .ip2(n17333), .s(n17410), .op(n17306) );
  mux2_1 U17365 ( .ip1(\x[119][14] ), .ip2(n17334), .s(n17410), .op(n17305) );
  mux2_1 U17366 ( .ip1(\x[119][13] ), .ip2(n17335), .s(n17410), .op(n17304) );
  mux2_1 U17367 ( .ip1(\x[119][12] ), .ip2(n17336), .s(n17410), .op(n17303) );
  mux2_1 U17368 ( .ip1(\x[119][11] ), .ip2(n17337), .s(n17410), .op(n17302) );
  mux2_1 U17369 ( .ip1(\x[119][10] ), .ip2(n17338), .s(n17410), .op(n17301) );
  buf_1 U17370 ( .ip(n17410), .op(n17409) );
  mux2_1 U17371 ( .ip1(\x[119][9] ), .ip2(n17339), .s(n17409), .op(n17300) );
  mux2_1 U17372 ( .ip1(\x[119][8] ), .ip2(n17340), .s(n17410), .op(n17299) );
  mux2_1 U17373 ( .ip1(\x[119][7] ), .ip2(n17341), .s(n17409), .op(n17298) );
  mux2_1 U17374 ( .ip1(\x[119][6] ), .ip2(n17342), .s(n17410), .op(n17297) );
  mux2_1 U17375 ( .ip1(\x[119][5] ), .ip2(n17343), .s(n17409), .op(n17296) );
  mux2_1 U17376 ( .ip1(\x[119][4] ), .ip2(n17344), .s(n17410), .op(n17295) );
  mux2_1 U17377 ( .ip1(\x[119][3] ), .ip2(n17345), .s(n17409), .op(n17294) );
  mux2_1 U17378 ( .ip1(\x[119][2] ), .ip2(n17346), .s(n17409), .op(n17293) );
  mux2_1 U17379 ( .ip1(\x[119][1] ), .ip2(n17347), .s(n17409), .op(n17292) );
  mux2_1 U17380 ( .ip1(\x[119][0] ), .ip2(n17348), .s(n17409), .op(n17291) );
  nor2_1 U17381 ( .ip1(address[0]), .ip2(address[3]), .op(n17325) );
  nand3_1 U17382 ( .ip1(address[2]), .ip2(address[1]), .ip3(n17325), .op(
        n17398) );
  nor2_1 U17383 ( .ip1(n17326), .ip2(n17398), .op(n17412) );
  mux2_1 U17384 ( .ip1(\x[118][15] ), .ip2(n17333), .s(n17412), .op(n17290) );
  mux2_1 U17385 ( .ip1(\x[118][14] ), .ip2(n17334), .s(n17412), .op(n17289) );
  mux2_1 U17386 ( .ip1(\x[118][13] ), .ip2(n17335), .s(n17412), .op(n17288) );
  mux2_1 U17387 ( .ip1(\x[118][12] ), .ip2(n17336), .s(n17412), .op(n17287) );
  mux2_1 U17388 ( .ip1(\x[118][11] ), .ip2(n17337), .s(n17412), .op(n17286) );
  mux2_1 U17389 ( .ip1(\x[118][10] ), .ip2(n17338), .s(n17412), .op(n17285) );
  buf_1 U17390 ( .ip(n17412), .op(n17411) );
  mux2_1 U17391 ( .ip1(\x[118][9] ), .ip2(n17339), .s(n17411), .op(n17284) );
  mux2_1 U17392 ( .ip1(\x[118][8] ), .ip2(n17340), .s(n17412), .op(n17283) );
  mux2_1 U17393 ( .ip1(\x[118][7] ), .ip2(n17341), .s(n17411), .op(n17282) );
  mux2_1 U17394 ( .ip1(\x[118][6] ), .ip2(n17342), .s(n17412), .op(n17281) );
  mux2_1 U17395 ( .ip1(\x[118][5] ), .ip2(n17343), .s(n17411), .op(n17280) );
  mux2_1 U17396 ( .ip1(\x[118][4] ), .ip2(n17344), .s(n17412), .op(n17279) );
  mux2_1 U17397 ( .ip1(\x[118][3] ), .ip2(n17345), .s(n17411), .op(n17278) );
  mux2_1 U17398 ( .ip1(\x[118][2] ), .ip2(n17346), .s(n17411), .op(n17277) );
  mux2_1 U17399 ( .ip1(\x[118][1] ), .ip2(n17347), .s(n17411), .op(n17276) );
  mux2_1 U17400 ( .ip1(\x[118][0] ), .ip2(n17348), .s(n17411), .op(n17275) );
  inv_1 U17401 ( .ip(address[2]), .op(n17329) );
  nor2_1 U17402 ( .ip1(address[1]), .ip2(n17329), .op(n17328) );
  nand3_1 U17403 ( .ip1(address[0]), .ip2(n17328), .ip3(n17324), .op(n17399)
         );
  nor2_1 U17404 ( .ip1(n17326), .ip2(n17399), .op(n17414) );
  mux2_1 U17405 ( .ip1(\x[117][15] ), .ip2(n17333), .s(n17414), .op(n17274) );
  mux2_1 U17406 ( .ip1(\x[117][14] ), .ip2(n17334), .s(n17414), .op(n17273) );
  mux2_1 U17407 ( .ip1(\x[117][13] ), .ip2(n17335), .s(n17414), .op(n17272) );
  mux2_1 U17408 ( .ip1(\x[117][12] ), .ip2(n17336), .s(n17414), .op(n17271) );
  mux2_1 U17409 ( .ip1(\x[117][11] ), .ip2(n17337), .s(n17414), .op(n17270) );
  mux2_1 U17410 ( .ip1(\x[117][10] ), .ip2(n17338), .s(n17414), .op(n17269) );
  buf_1 U17411 ( .ip(n17414), .op(n17413) );
  mux2_1 U17412 ( .ip1(\x[117][9] ), .ip2(n17339), .s(n17413), .op(n17268) );
  mux2_1 U17413 ( .ip1(\x[117][8] ), .ip2(n17340), .s(n17414), .op(n17267) );
  mux2_1 U17414 ( .ip1(\x[117][7] ), .ip2(n17341), .s(n17413), .op(n17266) );
  mux2_1 U17415 ( .ip1(\x[117][6] ), .ip2(n17342), .s(n17414), .op(n17265) );
  mux2_1 U17416 ( .ip1(\x[117][5] ), .ip2(n17343), .s(n17413), .op(n17264) );
  mux2_1 U17417 ( .ip1(\x[117][4] ), .ip2(n17344), .s(n17414), .op(n17263) );
  mux2_1 U17418 ( .ip1(\x[117][3] ), .ip2(n17345), .s(n17413), .op(n17262) );
  mux2_1 U17419 ( .ip1(\x[117][2] ), .ip2(n17346), .s(n17413), .op(n17261) );
  mux2_1 U17420 ( .ip1(\x[117][1] ), .ip2(n17347), .s(n17413), .op(n17260) );
  mux2_1 U17421 ( .ip1(\x[117][0] ), .ip2(n17348), .s(n17413), .op(n17259) );
  nand2_1 U17422 ( .ip1(n17325), .ip2(n17328), .op(n17400) );
  nor2_1 U17423 ( .ip1(n17326), .ip2(n17400), .op(n17416) );
  mux2_1 U17424 ( .ip1(\x[116][15] ), .ip2(n17333), .s(n17416), .op(n17258) );
  mux2_1 U17425 ( .ip1(\x[116][14] ), .ip2(n17334), .s(n17416), .op(n17257) );
  mux2_1 U17426 ( .ip1(\x[116][13] ), .ip2(n17335), .s(n17416), .op(n17256) );
  mux2_1 U17427 ( .ip1(\x[116][12] ), .ip2(n17336), .s(n17416), .op(n17255) );
  mux2_1 U17428 ( .ip1(\x[116][11] ), .ip2(n17337), .s(n17416), .op(n17254) );
  mux2_1 U17429 ( .ip1(\x[116][10] ), .ip2(n17338), .s(n17416), .op(n17253) );
  buf_1 U17430 ( .ip(n17416), .op(n17415) );
  mux2_1 U17431 ( .ip1(\x[116][9] ), .ip2(n17339), .s(n17415), .op(n17252) );
  mux2_1 U17432 ( .ip1(\x[116][8] ), .ip2(n17340), .s(n17416), .op(n17251) );
  mux2_1 U17433 ( .ip1(\x[116][7] ), .ip2(n17341), .s(n17415), .op(n17250) );
  mux2_1 U17434 ( .ip1(\x[116][6] ), .ip2(n17342), .s(n17416), .op(n17249) );
  mux2_1 U17435 ( .ip1(\x[116][5] ), .ip2(n17343), .s(n17415), .op(n17248) );
  mux2_1 U17436 ( .ip1(\x[116][4] ), .ip2(n17344), .s(n17416), .op(n17247) );
  mux2_1 U17437 ( .ip1(\x[116][3] ), .ip2(n17345), .s(n17415), .op(n17246) );
  mux2_1 U17438 ( .ip1(\x[116][2] ), .ip2(n17346), .s(n17415), .op(n17245) );
  mux2_1 U17439 ( .ip1(\x[116][1] ), .ip2(n17347), .s(n17415), .op(n17244) );
  mux2_1 U17440 ( .ip1(\x[116][0] ), .ip2(n17348), .s(n17415), .op(n17243) );
  nand4_1 U17441 ( .ip1(address[1]), .ip2(address[0]), .ip3(n17329), .ip4(
        n17324), .op(n17401) );
  nor2_1 U17442 ( .ip1(n17326), .ip2(n17401), .op(n17418) );
  mux2_1 U17443 ( .ip1(\x[115][15] ), .ip2(n17333), .s(n17418), .op(n17242) );
  mux2_1 U17444 ( .ip1(\x[115][14] ), .ip2(n17334), .s(n17418), .op(n17241) );
  mux2_1 U17445 ( .ip1(\x[115][13] ), .ip2(n17335), .s(n17418), .op(n17240) );
  mux2_1 U17446 ( .ip1(\x[115][12] ), .ip2(n17336), .s(n17418), .op(n17239) );
  mux2_1 U17447 ( .ip1(\x[115][11] ), .ip2(n17337), .s(n17418), .op(n17238) );
  mux2_1 U17448 ( .ip1(\x[115][10] ), .ip2(n17338), .s(n17418), .op(n17237) );
  buf_1 U17449 ( .ip(n17418), .op(n17417) );
  mux2_1 U17450 ( .ip1(\x[115][9] ), .ip2(n17339), .s(n17417), .op(n17236) );
  mux2_1 U17451 ( .ip1(\x[115][8] ), .ip2(n17340), .s(n17418), .op(n17235) );
  mux2_1 U17452 ( .ip1(\x[115][7] ), .ip2(n17341), .s(n17417), .op(n17234) );
  mux2_1 U17453 ( .ip1(\x[115][6] ), .ip2(n17342), .s(n17418), .op(n17233) );
  mux2_1 U17454 ( .ip1(\x[115][5] ), .ip2(n17343), .s(n17417), .op(n17232) );
  mux2_1 U17455 ( .ip1(\x[115][4] ), .ip2(n17344), .s(n17418), .op(n17231) );
  mux2_1 U17456 ( .ip1(\x[115][3] ), .ip2(n17345), .s(n17417), .op(n17230) );
  mux2_1 U17457 ( .ip1(\x[115][2] ), .ip2(n17346), .s(n17417), .op(n17229) );
  mux2_1 U17458 ( .ip1(\x[115][1] ), .ip2(n17347), .s(n17417), .op(n17228) );
  mux2_1 U17459 ( .ip1(\x[115][0] ), .ip2(n17348), .s(n17417), .op(n17227) );
  nand3_1 U17460 ( .ip1(address[1]), .ip2(n17325), .ip3(n17329), .op(n17402)
         );
  nor2_1 U17461 ( .ip1(n17326), .ip2(n17402), .op(n17420) );
  mux2_1 U17462 ( .ip1(\x[114][15] ), .ip2(n17333), .s(n17420), .op(n17226) );
  mux2_1 U17463 ( .ip1(\x[114][14] ), .ip2(n17334), .s(n17420), .op(n17225) );
  mux2_1 U17464 ( .ip1(\x[114][13] ), .ip2(n17335), .s(n17420), .op(n17224) );
  mux2_1 U17465 ( .ip1(\x[114][12] ), .ip2(n17336), .s(n17420), .op(n17223) );
  mux2_1 U17466 ( .ip1(\x[114][11] ), .ip2(n17337), .s(n17420), .op(n17222) );
  mux2_1 U17467 ( .ip1(\x[114][10] ), .ip2(n17338), .s(n17420), .op(n17221) );
  buf_1 U17468 ( .ip(n17420), .op(n17419) );
  mux2_1 U17469 ( .ip1(\x[114][9] ), .ip2(n17339), .s(n17419), .op(n17220) );
  mux2_1 U17470 ( .ip1(\x[114][8] ), .ip2(n17340), .s(n17420), .op(n17219) );
  mux2_1 U17471 ( .ip1(\x[114][7] ), .ip2(n17341), .s(n17419), .op(n17218) );
  mux2_1 U17472 ( .ip1(\x[114][6] ), .ip2(n17342), .s(n17420), .op(n17217) );
  mux2_1 U17473 ( .ip1(\x[114][5] ), .ip2(n17343), .s(n17419), .op(n17216) );
  mux2_1 U17474 ( .ip1(\x[114][4] ), .ip2(n17344), .s(n17420), .op(n17215) );
  mux2_1 U17475 ( .ip1(\x[114][3] ), .ip2(n17345), .s(n17419), .op(n17214) );
  mux2_1 U17476 ( .ip1(\x[114][2] ), .ip2(n17346), .s(n17419), .op(n17213) );
  mux2_1 U17477 ( .ip1(\x[114][1] ), .ip2(n17347), .s(n17419), .op(n17212) );
  mux2_1 U17478 ( .ip1(\x[114][0] ), .ip2(n17348), .s(n17419), .op(n17211) );
  nand3_1 U17479 ( .ip1(address[0]), .ip2(n17331), .ip3(n17324), .op(n17403)
         );
  nor2_1 U17480 ( .ip1(n17326), .ip2(n17403), .op(n17422) );
  mux2_1 U17481 ( .ip1(\x[113][15] ), .ip2(n17333), .s(n17422), .op(n17210) );
  mux2_1 U17482 ( .ip1(\x[113][14] ), .ip2(n17334), .s(n17422), .op(n17209) );
  mux2_1 U17483 ( .ip1(\x[113][13] ), .ip2(n17335), .s(n17422), .op(n17208) );
  mux2_1 U17484 ( .ip1(\x[113][12] ), .ip2(n17336), .s(n17422), .op(n17207) );
  mux2_1 U17485 ( .ip1(\x[113][11] ), .ip2(n17337), .s(n17422), .op(n17206) );
  mux2_1 U17486 ( .ip1(\x[113][10] ), .ip2(n17338), .s(n17422), .op(n17205) );
  buf_1 U17487 ( .ip(n17422), .op(n17421) );
  mux2_1 U17488 ( .ip1(\x[113][9] ), .ip2(n17339), .s(n17421), .op(n17204) );
  mux2_1 U17489 ( .ip1(\x[113][8] ), .ip2(n17340), .s(n17422), .op(n17203) );
  mux2_1 U17490 ( .ip1(\x[113][7] ), .ip2(n17341), .s(n17421), .op(n17202) );
  mux2_1 U17491 ( .ip1(\x[113][6] ), .ip2(n17342), .s(n17422), .op(n17201) );
  mux2_1 U17492 ( .ip1(\x[113][5] ), .ip2(n17343), .s(n17421), .op(n17200) );
  mux2_1 U17493 ( .ip1(\x[113][4] ), .ip2(n17344), .s(n17422), .op(n17199) );
  mux2_1 U17494 ( .ip1(\x[113][3] ), .ip2(n17345), .s(n17421), .op(n17198) );
  mux2_1 U17495 ( .ip1(\x[113][2] ), .ip2(n17346), .s(n17421), .op(n17197) );
  mux2_1 U17496 ( .ip1(\x[113][1] ), .ip2(n17347), .s(n17421), .op(n17196) );
  mux2_1 U17497 ( .ip1(\x[113][0] ), .ip2(n17348), .s(n17421), .op(n17195) );
  nand2_1 U17498 ( .ip1(n17331), .ip2(n17325), .op(n17405) );
  nor2_1 U17499 ( .ip1(n17326), .ip2(n17405), .op(n17424) );
  mux2_1 U17500 ( .ip1(\x[112][15] ), .ip2(n17333), .s(n17424), .op(n17194) );
  mux2_1 U17501 ( .ip1(\x[112][14] ), .ip2(n17334), .s(n17424), .op(n17193) );
  mux2_1 U17502 ( .ip1(\x[112][13] ), .ip2(n17335), .s(n17424), .op(n17192) );
  mux2_1 U17503 ( .ip1(\x[112][12] ), .ip2(n17336), .s(n17424), .op(n17191) );
  mux2_1 U17504 ( .ip1(\x[112][11] ), .ip2(n17337), .s(n17424), .op(n17190) );
  mux2_1 U17505 ( .ip1(\x[112][10] ), .ip2(n17338), .s(n17424), .op(n17189) );
  buf_1 U17506 ( .ip(n17424), .op(n17423) );
  mux2_1 U17507 ( .ip1(\x[112][9] ), .ip2(n17339), .s(n17423), .op(n17188) );
  mux2_1 U17508 ( .ip1(\x[112][8] ), .ip2(n17340), .s(n17424), .op(n17187) );
  mux2_1 U17509 ( .ip1(\x[112][7] ), .ip2(n17341), .s(n17423), .op(n17186) );
  mux2_1 U17510 ( .ip1(\x[112][6] ), .ip2(n17342), .s(n17424), .op(n17185) );
  mux2_1 U17511 ( .ip1(\x[112][5] ), .ip2(n17343), .s(n17423), .op(n17184) );
  mux2_1 U17512 ( .ip1(\x[112][4] ), .ip2(n17344), .s(n17424), .op(n17183) );
  mux2_1 U17513 ( .ip1(\x[112][3] ), .ip2(n17345), .s(n17423), .op(n17182) );
  mux2_1 U17514 ( .ip1(\x[112][2] ), .ip2(n17346), .s(n17423), .op(n17181) );
  mux2_1 U17515 ( .ip1(\x[112][1] ), .ip2(n17347), .s(n17423), .op(n17180) );
  mux2_1 U17516 ( .ip1(\x[112][0] ), .ip2(n17348), .s(n17423), .op(n17179) );
  nand4_1 U17517 ( .ip1(address[2]), .ip2(address[1]), .ip3(address[0]), .ip4(
        address[3]), .op(n17373) );
  inv_1 U17518 ( .ip(we), .op(n17327) );
  nor2_1 U17519 ( .ip1(address[4]), .ip2(n17327), .op(n17372) );
  nand3_1 U17520 ( .ip1(address[6]), .ip2(address[5]), .ip3(n17372), .op(
        n17332) );
  nor2_1 U17521 ( .ip1(n17373), .ip2(n17332), .op(n17426) );
  mux2_1 U17522 ( .ip1(\x[111][15] ), .ip2(n17333), .s(n17426), .op(n17178) );
  mux2_1 U17523 ( .ip1(\x[111][14] ), .ip2(n17334), .s(n17426), .op(n17177) );
  mux2_1 U17524 ( .ip1(\x[111][13] ), .ip2(n17335), .s(n17426), .op(n17176) );
  mux2_1 U17525 ( .ip1(\x[111][12] ), .ip2(n17336), .s(n17426), .op(n17175) );
  mux2_1 U17526 ( .ip1(\x[111][11] ), .ip2(n17337), .s(n17426), .op(n17174) );
  mux2_1 U17527 ( .ip1(\x[111][10] ), .ip2(n17338), .s(n17426), .op(n17173) );
  buf_1 U17528 ( .ip(n17426), .op(n17425) );
  mux2_1 U17529 ( .ip1(\x[111][9] ), .ip2(n17339), .s(n17425), .op(n17172) );
  mux2_1 U17530 ( .ip1(\x[111][8] ), .ip2(n17340), .s(n17426), .op(n17171) );
  mux2_1 U17531 ( .ip1(\x[111][7] ), .ip2(n17341), .s(n17425), .op(n17170) );
  mux2_1 U17532 ( .ip1(\x[111][6] ), .ip2(n17342), .s(n17426), .op(n17169) );
  mux2_1 U17533 ( .ip1(\x[111][5] ), .ip2(n17343), .s(n17425), .op(n17168) );
  mux2_1 U17534 ( .ip1(\x[111][4] ), .ip2(n17344), .s(n17426), .op(n17167) );
  mux2_1 U17535 ( .ip1(\x[111][3] ), .ip2(n17345), .s(n17425), .op(n17166) );
  mux2_1 U17536 ( .ip1(\x[111][2] ), .ip2(n17346), .s(n17425), .op(n17165) );
  mux2_1 U17537 ( .ip1(\x[111][1] ), .ip2(n17347), .s(n17425), .op(n17164) );
  mux2_1 U17538 ( .ip1(\x[111][0] ), .ip2(n17348), .s(n17425), .op(n17163) );
  nand3_1 U17539 ( .ip1(address[2]), .ip2(address[1]), .ip3(n17330), .op(
        n17374) );
  nor2_1 U17540 ( .ip1(n17332), .ip2(n17374), .op(n17428) );
  mux2_1 U17541 ( .ip1(\x[110][15] ), .ip2(n17333), .s(n17428), .op(n17162) );
  mux2_1 U17542 ( .ip1(\x[110][14] ), .ip2(n17334), .s(n17428), .op(n17161) );
  mux2_1 U17543 ( .ip1(\x[110][13] ), .ip2(n17335), .s(n17428), .op(n17160) );
  mux2_1 U17544 ( .ip1(\x[110][12] ), .ip2(n17336), .s(n17428), .op(n17159) );
  mux2_1 U17545 ( .ip1(\x[110][11] ), .ip2(n17337), .s(n17428), .op(n17158) );
  mux2_1 U17546 ( .ip1(\x[110][10] ), .ip2(n17338), .s(n17428), .op(n17157) );
  buf_1 U17547 ( .ip(n17428), .op(n17427) );
  mux2_1 U17548 ( .ip1(\x[110][9] ), .ip2(n17339), .s(n17427), .op(n17156) );
  mux2_1 U17549 ( .ip1(\x[110][8] ), .ip2(n17340), .s(n17428), .op(n17155) );
  mux2_1 U17550 ( .ip1(\x[110][7] ), .ip2(n17341), .s(n17427), .op(n17154) );
  mux2_1 U17551 ( .ip1(\x[110][6] ), .ip2(n17342), .s(n17428), .op(n17153) );
  mux2_1 U17552 ( .ip1(\x[110][5] ), .ip2(n17343), .s(n17427), .op(n17152) );
  mux2_1 U17553 ( .ip1(\x[110][4] ), .ip2(n17344), .s(n17428), .op(n17151) );
  mux2_1 U17554 ( .ip1(\x[110][3] ), .ip2(n17345), .s(n17427), .op(n17150) );
  mux2_1 U17555 ( .ip1(\x[110][2] ), .ip2(n17346), .s(n17427), .op(n17149) );
  mux2_1 U17556 ( .ip1(\x[110][1] ), .ip2(n17347), .s(n17427), .op(n17148) );
  mux2_1 U17557 ( .ip1(\x[110][0] ), .ip2(n17348), .s(n17427), .op(n17147) );
  nand3_1 U17558 ( .ip1(address[0]), .ip2(address[3]), .ip3(n17328), .op(
        n17375) );
  nor2_1 U17559 ( .ip1(n17332), .ip2(n17375), .op(n17430) );
  mux2_1 U17560 ( .ip1(\x[109][15] ), .ip2(n17333), .s(n17430), .op(n17146) );
  mux2_1 U17561 ( .ip1(\x[109][14] ), .ip2(n17334), .s(n17430), .op(n17145) );
  mux2_1 U17562 ( .ip1(\x[109][13] ), .ip2(n17335), .s(n17430), .op(n17144) );
  mux2_1 U17563 ( .ip1(\x[109][12] ), .ip2(n17336), .s(n17430), .op(n17143) );
  mux2_1 U17564 ( .ip1(\x[109][11] ), .ip2(n17337), .s(n17430), .op(n17142) );
  mux2_1 U17565 ( .ip1(\x[109][10] ), .ip2(n17338), .s(n17430), .op(n17141) );
  buf_1 U17566 ( .ip(n17430), .op(n17429) );
  mux2_1 U17567 ( .ip1(\x[109][9] ), .ip2(n17339), .s(n17429), .op(n17140) );
  mux2_1 U17568 ( .ip1(\x[109][8] ), .ip2(n17340), .s(n17430), .op(n17139) );
  mux2_1 U17569 ( .ip1(\x[109][7] ), .ip2(n17341), .s(n17429), .op(n17138) );
  mux2_1 U17570 ( .ip1(\x[109][6] ), .ip2(n17342), .s(n17430), .op(n17137) );
  mux2_1 U17571 ( .ip1(\x[109][5] ), .ip2(n17343), .s(n17429), .op(n17136) );
  mux2_1 U17572 ( .ip1(\x[109][4] ), .ip2(n17344), .s(n17430), .op(n17135) );
  mux2_1 U17573 ( .ip1(\x[109][3] ), .ip2(n17345), .s(n17429), .op(n17134) );
  mux2_1 U17574 ( .ip1(\x[109][2] ), .ip2(n17346), .s(n17429), .op(n17133) );
  mux2_1 U17575 ( .ip1(\x[109][1] ), .ip2(n17347), .s(n17429), .op(n17132) );
  mux2_1 U17576 ( .ip1(\x[109][0] ), .ip2(n17348), .s(n17429), .op(n17131) );
  nand2_1 U17577 ( .ip1(n17330), .ip2(n17328), .op(n17392) );
  nor2_1 U17578 ( .ip1(n17332), .ip2(n17392), .op(n17432) );
  mux2_1 U17579 ( .ip1(\x[108][15] ), .ip2(n17333), .s(n17432), .op(n17130) );
  mux2_1 U17580 ( .ip1(\x[108][14] ), .ip2(n17334), .s(n17432), .op(n17129) );
  mux2_1 U17581 ( .ip1(\x[108][13] ), .ip2(n17335), .s(n17432), .op(n17128) );
  mux2_1 U17582 ( .ip1(\x[108][12] ), .ip2(n17336), .s(n17432), .op(n17127) );
  mux2_1 U17583 ( .ip1(\x[108][11] ), .ip2(n17337), .s(n17432), .op(n17126) );
  mux2_1 U17584 ( .ip1(\x[108][10] ), .ip2(n17338), .s(n17432), .op(n17125) );
  buf_1 U17585 ( .ip(n17432), .op(n17431) );
  mux2_1 U17586 ( .ip1(\x[108][9] ), .ip2(n17339), .s(n17431), .op(n17124) );
  mux2_1 U17587 ( .ip1(\x[108][8] ), .ip2(n17340), .s(n17432), .op(n17123) );
  mux2_1 U17588 ( .ip1(\x[108][7] ), .ip2(n17341), .s(n17431), .op(n17122) );
  mux2_1 U17589 ( .ip1(\x[108][6] ), .ip2(n17342), .s(n17432), .op(n17121) );
  mux2_1 U17590 ( .ip1(\x[108][5] ), .ip2(n17343), .s(n17431), .op(n17120) );
  mux2_1 U17591 ( .ip1(\x[108][4] ), .ip2(n17344), .s(n17432), .op(n17119) );
  mux2_1 U17592 ( .ip1(\x[108][3] ), .ip2(n17345), .s(n17431), .op(n17118) );
  mux2_1 U17593 ( .ip1(\x[108][2] ), .ip2(n17346), .s(n17431), .op(n17117) );
  mux2_1 U17594 ( .ip1(\x[108][1] ), .ip2(n17347), .s(n17431), .op(n17116) );
  mux2_1 U17595 ( .ip1(\x[108][0] ), .ip2(n17348), .s(n17431), .op(n17115) );
  nand4_1 U17596 ( .ip1(address[1]), .ip2(address[0]), .ip3(address[3]), .ip4(
        n17329), .op(n17393) );
  nor2_1 U17597 ( .ip1(n17332), .ip2(n17393), .op(n17434) );
  mux2_1 U17598 ( .ip1(\x[107][15] ), .ip2(n17333), .s(n17434), .op(n17114) );
  mux2_1 U17599 ( .ip1(\x[107][14] ), .ip2(n17334), .s(n17434), .op(n17113) );
  mux2_1 U17600 ( .ip1(\x[107][13] ), .ip2(n17335), .s(n17434), .op(n17112) );
  mux2_1 U17601 ( .ip1(\x[107][12] ), .ip2(n17336), .s(n17434), .op(n17111) );
  mux2_1 U17602 ( .ip1(\x[107][11] ), .ip2(n17337), .s(n17434), .op(n17110) );
  mux2_1 U17603 ( .ip1(\x[107][10] ), .ip2(n17338), .s(n17434), .op(n17109) );
  buf_1 U17604 ( .ip(n17434), .op(n17433) );
  mux2_1 U17605 ( .ip1(\x[107][9] ), .ip2(n17339), .s(n17433), .op(n17108) );
  mux2_1 U17606 ( .ip1(\x[107][8] ), .ip2(n17340), .s(n17434), .op(n17107) );
  mux2_1 U17607 ( .ip1(\x[107][7] ), .ip2(n17341), .s(n17433), .op(n17106) );
  mux2_1 U17608 ( .ip1(\x[107][6] ), .ip2(n17342), .s(n17434), .op(n17105) );
  mux2_1 U17609 ( .ip1(\x[107][5] ), .ip2(n17343), .s(n17433), .op(n17104) );
  mux2_1 U17610 ( .ip1(\x[107][4] ), .ip2(n17344), .s(n17434), .op(n17103) );
  mux2_1 U17611 ( .ip1(\x[107][3] ), .ip2(n17345), .s(n17433), .op(n17102) );
  mux2_1 U17612 ( .ip1(\x[107][2] ), .ip2(n17346), .s(n17433), .op(n17101) );
  mux2_1 U17613 ( .ip1(\x[107][1] ), .ip2(n17347), .s(n17433), .op(n17100) );
  mux2_1 U17614 ( .ip1(\x[107][0] ), .ip2(n17348), .s(n17433), .op(n17099) );
  nand3_1 U17615 ( .ip1(address[1]), .ip2(n17330), .ip3(n17329), .op(n17394)
         );
  nor2_1 U17616 ( .ip1(n17332), .ip2(n17394), .op(n17436) );
  mux2_1 U17617 ( .ip1(\x[106][15] ), .ip2(n17333), .s(n17436), .op(n17098) );
  mux2_1 U17618 ( .ip1(\x[106][14] ), .ip2(n17334), .s(n17436), .op(n17097) );
  mux2_1 U17619 ( .ip1(\x[106][13] ), .ip2(n17335), .s(n17436), .op(n17096) );
  mux2_1 U17620 ( .ip1(\x[106][12] ), .ip2(n17336), .s(n17436), .op(n17095) );
  mux2_1 U17621 ( .ip1(\x[106][11] ), .ip2(n17337), .s(n17436), .op(n17094) );
  mux2_1 U17622 ( .ip1(\x[106][10] ), .ip2(n17338), .s(n17436), .op(n17093) );
  buf_1 U17623 ( .ip(n17436), .op(n17435) );
  mux2_1 U17624 ( .ip1(\x[106][9] ), .ip2(n17339), .s(n17435), .op(n17092) );
  mux2_1 U17625 ( .ip1(\x[106][8] ), .ip2(n17340), .s(n17436), .op(n17091) );
  mux2_1 U17626 ( .ip1(\x[106][7] ), .ip2(n17341), .s(n17435), .op(n17090) );
  mux2_1 U17627 ( .ip1(\x[106][6] ), .ip2(n17342), .s(n17436), .op(n17089) );
  mux2_1 U17628 ( .ip1(\x[106][5] ), .ip2(n17343), .s(n17435), .op(n17088) );
  mux2_1 U17629 ( .ip1(\x[106][4] ), .ip2(n17344), .s(n17436), .op(n17087) );
  mux2_1 U17630 ( .ip1(\x[106][3] ), .ip2(n17345), .s(n17435), .op(n17086) );
  mux2_1 U17631 ( .ip1(\x[106][2] ), .ip2(n17346), .s(n17435), .op(n17085) );
  mux2_1 U17632 ( .ip1(\x[106][1] ), .ip2(n17347), .s(n17435), .op(n17084) );
  mux2_1 U17633 ( .ip1(\x[106][0] ), .ip2(n17348), .s(n17435), .op(n17083) );
  nand3_1 U17634 ( .ip1(n17331), .ip2(address[0]), .ip3(address[3]), .op(
        n17395) );
  nor2_1 U17635 ( .ip1(n17332), .ip2(n17395), .op(n17438) );
  mux2_1 U17636 ( .ip1(\x[105][15] ), .ip2(n17333), .s(n17438), .op(n17082) );
  mux2_1 U17637 ( .ip1(\x[105][14] ), .ip2(n17334), .s(n17438), .op(n17081) );
  mux2_1 U17638 ( .ip1(\x[105][13] ), .ip2(n17335), .s(n17438), .op(n17080) );
  mux2_1 U17639 ( .ip1(\x[105][12] ), .ip2(n17336), .s(n17438), .op(n17079) );
  mux2_1 U17640 ( .ip1(\x[105][11] ), .ip2(n17337), .s(n17438), .op(n17078) );
  mux2_1 U17641 ( .ip1(\x[105][10] ), .ip2(n17338), .s(n17438), .op(n17077) );
  buf_1 U17642 ( .ip(n17438), .op(n17437) );
  mux2_1 U17643 ( .ip1(\x[105][9] ), .ip2(n17339), .s(n17437), .op(n17076) );
  mux2_1 U17644 ( .ip1(\x[105][8] ), .ip2(n17340), .s(n17438), .op(n17075) );
  mux2_1 U17645 ( .ip1(\x[105][7] ), .ip2(n17341), .s(n17437), .op(n17074) );
  mux2_1 U17646 ( .ip1(\x[105][6] ), .ip2(n17342), .s(n17438), .op(n17073) );
  mux2_1 U17647 ( .ip1(\x[105][5] ), .ip2(n17343), .s(n17437), .op(n17072) );
  mux2_1 U17648 ( .ip1(\x[105][4] ), .ip2(n17344), .s(n17438), .op(n17071) );
  mux2_1 U17649 ( .ip1(\x[105][3] ), .ip2(n17345), .s(n17437), .op(n17070) );
  mux2_1 U17650 ( .ip1(\x[105][2] ), .ip2(n17346), .s(n17437), .op(n17069) );
  mux2_1 U17651 ( .ip1(\x[105][1] ), .ip2(n17347), .s(n17437), .op(n17068) );
  mux2_1 U17652 ( .ip1(\x[105][0] ), .ip2(n17348), .s(n17437), .op(n17067) );
  nor2_1 U17653 ( .ip1(n17396), .ip2(n17332), .op(n17440) );
  mux2_1 U17654 ( .ip1(\x[104][15] ), .ip2(n17333), .s(n17440), .op(n17066) );
  mux2_1 U17655 ( .ip1(\x[104][14] ), .ip2(n17334), .s(n17440), .op(n17065) );
  mux2_1 U17656 ( .ip1(\x[104][13] ), .ip2(n17335), .s(n17440), .op(n17064) );
  mux2_1 U17657 ( .ip1(\x[104][12] ), .ip2(n17336), .s(n17440), .op(n17063) );
  mux2_1 U17658 ( .ip1(\x[104][11] ), .ip2(n17337), .s(n17440), .op(n17062) );
  mux2_1 U17659 ( .ip1(\x[104][10] ), .ip2(n17338), .s(n17440), .op(n17061) );
  buf_1 U17660 ( .ip(n17440), .op(n17439) );
  mux2_1 U17661 ( .ip1(\x[104][9] ), .ip2(n17339), .s(n17439), .op(n17060) );
  mux2_1 U17662 ( .ip1(\x[104][8] ), .ip2(n17340), .s(n17440), .op(n17059) );
  mux2_1 U17663 ( .ip1(\x[104][7] ), .ip2(n17341), .s(n17439), .op(n17058) );
  mux2_1 U17664 ( .ip1(\x[104][6] ), .ip2(n17342), .s(n17440), .op(n17057) );
  mux2_1 U17665 ( .ip1(\x[104][5] ), .ip2(n17343), .s(n17439), .op(n17056) );
  mux2_1 U17666 ( .ip1(\x[104][4] ), .ip2(n17344), .s(n17440), .op(n17055) );
  mux2_1 U17667 ( .ip1(\x[104][3] ), .ip2(n17345), .s(n17439), .op(n17054) );
  mux2_1 U17668 ( .ip1(\x[104][2] ), .ip2(n17346), .s(n17439), .op(n17053) );
  mux2_1 U17669 ( .ip1(\x[104][1] ), .ip2(n17347), .s(n17439), .op(n17052) );
  mux2_1 U17670 ( .ip1(\x[104][0] ), .ip2(n17348), .s(n17439), .op(n17051) );
  nor2_1 U17671 ( .ip1(n17397), .ip2(n17332), .op(n17442) );
  mux2_1 U17672 ( .ip1(\x[103][15] ), .ip2(n17333), .s(n17442), .op(n17050) );
  mux2_1 U17673 ( .ip1(\x[103][14] ), .ip2(n17334), .s(n17442), .op(n17049) );
  mux2_1 U17674 ( .ip1(\x[103][13] ), .ip2(n17335), .s(n17442), .op(n17048) );
  mux2_1 U17675 ( .ip1(\x[103][12] ), .ip2(n17336), .s(n17442), .op(n17047) );
  mux2_1 U17676 ( .ip1(\x[103][11] ), .ip2(n17337), .s(n17442), .op(n17046) );
  mux2_1 U17677 ( .ip1(\x[103][10] ), .ip2(n17338), .s(n17442), .op(n17045) );
  buf_1 U17678 ( .ip(n17442), .op(n17441) );
  mux2_1 U17679 ( .ip1(\x[103][9] ), .ip2(n17339), .s(n17441), .op(n17044) );
  mux2_1 U17680 ( .ip1(\x[103][8] ), .ip2(n17340), .s(n17442), .op(n17043) );
  mux2_1 U17681 ( .ip1(\x[103][7] ), .ip2(n17341), .s(n17441), .op(n17042) );
  mux2_1 U17682 ( .ip1(\x[103][6] ), .ip2(n17342), .s(n17442), .op(n17041) );
  mux2_1 U17683 ( .ip1(\x[103][5] ), .ip2(n17343), .s(n17441), .op(n17040) );
  mux2_1 U17684 ( .ip1(\x[103][4] ), .ip2(n17344), .s(n17442), .op(n17039) );
  mux2_1 U17685 ( .ip1(\x[103][3] ), .ip2(n17345), .s(n17441), .op(n17038) );
  mux2_1 U17686 ( .ip1(\x[103][2] ), .ip2(n17346), .s(n17441), .op(n17037) );
  mux2_1 U17687 ( .ip1(\x[103][1] ), .ip2(n17347), .s(n17441), .op(n17036) );
  mux2_1 U17688 ( .ip1(\x[103][0] ), .ip2(n17348), .s(n17441), .op(n17035) );
  nor2_1 U17689 ( .ip1(n17398), .ip2(n17332), .op(n17444) );
  mux2_1 U17690 ( .ip1(\x[102][15] ), .ip2(n17333), .s(n17444), .op(n17034) );
  mux2_1 U17691 ( .ip1(\x[102][14] ), .ip2(n17334), .s(n17444), .op(n17033) );
  mux2_1 U17692 ( .ip1(\x[102][13] ), .ip2(n17335), .s(n17444), .op(n17032) );
  mux2_1 U17693 ( .ip1(\x[102][12] ), .ip2(n17336), .s(n17444), .op(n17031) );
  mux2_1 U17694 ( .ip1(\x[102][11] ), .ip2(n17337), .s(n17444), .op(n17030) );
  mux2_1 U17695 ( .ip1(\x[102][10] ), .ip2(n17338), .s(n17444), .op(n17029) );
  buf_1 U17696 ( .ip(n17444), .op(n17443) );
  mux2_1 U17697 ( .ip1(\x[102][9] ), .ip2(n17339), .s(n17443), .op(n17028) );
  mux2_1 U17698 ( .ip1(\x[102][8] ), .ip2(n17340), .s(n17444), .op(n17027) );
  mux2_1 U17699 ( .ip1(\x[102][7] ), .ip2(n17341), .s(n17443), .op(n17026) );
  mux2_1 U17700 ( .ip1(\x[102][6] ), .ip2(n17342), .s(n17444), .op(n17025) );
  mux2_1 U17701 ( .ip1(\x[102][5] ), .ip2(n17343), .s(n17443), .op(n17024) );
  mux2_1 U17702 ( .ip1(\x[102][4] ), .ip2(n17344), .s(n17444), .op(n17023) );
  mux2_1 U17703 ( .ip1(\x[102][3] ), .ip2(n17345), .s(n17443), .op(n17022) );
  mux2_1 U17704 ( .ip1(\x[102][2] ), .ip2(n17346), .s(n17443), .op(n17021) );
  mux2_1 U17705 ( .ip1(\x[102][1] ), .ip2(n17347), .s(n17443), .op(n17020) );
  mux2_1 U17706 ( .ip1(\x[102][0] ), .ip2(n17348), .s(n17443), .op(n17019) );
  nor2_1 U17707 ( .ip1(n17399), .ip2(n17332), .op(n17446) );
  mux2_1 U17708 ( .ip1(\x[101][15] ), .ip2(n17333), .s(n17446), .op(n17018) );
  mux2_1 U17709 ( .ip1(\x[101][14] ), .ip2(n17334), .s(n17446), .op(n17017) );
  mux2_1 U17710 ( .ip1(\x[101][13] ), .ip2(n17335), .s(n17446), .op(n17016) );
  mux2_1 U17711 ( .ip1(\x[101][12] ), .ip2(n17336), .s(n17446), .op(n17015) );
  mux2_1 U17712 ( .ip1(\x[101][11] ), .ip2(n17337), .s(n17446), .op(n17014) );
  mux2_1 U17713 ( .ip1(\x[101][10] ), .ip2(n17338), .s(n17446), .op(n17013) );
  buf_1 U17714 ( .ip(n17446), .op(n17445) );
  mux2_1 U17715 ( .ip1(\x[101][9] ), .ip2(n17339), .s(n17445), .op(n17012) );
  mux2_1 U17716 ( .ip1(\x[101][8] ), .ip2(n17340), .s(n17446), .op(n17011) );
  mux2_1 U17717 ( .ip1(\x[101][7] ), .ip2(n17341), .s(n17445), .op(n17010) );
  mux2_1 U17718 ( .ip1(\x[101][6] ), .ip2(n17342), .s(n17446), .op(n17009) );
  mux2_1 U17719 ( .ip1(\x[101][5] ), .ip2(n17343), .s(n17445), .op(n17008) );
  mux2_1 U17720 ( .ip1(\x[101][4] ), .ip2(n17344), .s(n17446), .op(n17007) );
  mux2_1 U17721 ( .ip1(\x[101][3] ), .ip2(n17345), .s(n17445), .op(n17006) );
  mux2_1 U17722 ( .ip1(\x[101][2] ), .ip2(n17346), .s(n17445), .op(n17005) );
  mux2_1 U17723 ( .ip1(\x[101][1] ), .ip2(n17347), .s(n17445), .op(n17004) );
  mux2_1 U17724 ( .ip1(\x[101][0] ), .ip2(n17348), .s(n17445), .op(n17003) );
  nor2_1 U17725 ( .ip1(n17400), .ip2(n17332), .op(n17448) );
  mux2_1 U17726 ( .ip1(\x[100][15] ), .ip2(n17333), .s(n17448), .op(n17002) );
  mux2_1 U17727 ( .ip1(\x[100][14] ), .ip2(n17334), .s(n17448), .op(n17001) );
  mux2_1 U17728 ( .ip1(\x[100][13] ), .ip2(n17335), .s(n17448), .op(n17000) );
  mux2_1 U17729 ( .ip1(\x[100][12] ), .ip2(n17336), .s(n17448), .op(n16999) );
  mux2_1 U17730 ( .ip1(\x[100][11] ), .ip2(n17337), .s(n17448), .op(n16998) );
  mux2_1 U17731 ( .ip1(\x[100][10] ), .ip2(n17338), .s(n17448), .op(n16997) );
  buf_1 U17732 ( .ip(n17448), .op(n17447) );
  mux2_1 U17733 ( .ip1(\x[100][9] ), .ip2(n17339), .s(n17447), .op(n16996) );
  mux2_1 U17734 ( .ip1(\x[100][8] ), .ip2(n17340), .s(n17448), .op(n16995) );
  mux2_1 U17735 ( .ip1(\x[100][7] ), .ip2(n17341), .s(n17447), .op(n16994) );
  mux2_1 U17736 ( .ip1(\x[100][6] ), .ip2(n17342), .s(n17448), .op(n16993) );
  mux2_1 U17737 ( .ip1(\x[100][5] ), .ip2(n17343), .s(n17447), .op(n16992) );
  mux2_1 U17738 ( .ip1(\x[100][4] ), .ip2(n17344), .s(n17448), .op(n16991) );
  mux2_1 U17739 ( .ip1(\x[100][3] ), .ip2(n17345), .s(n17447), .op(n16990) );
  mux2_1 U17740 ( .ip1(\x[100][2] ), .ip2(n17346), .s(n17447), .op(n16989) );
  mux2_1 U17741 ( .ip1(\x[100][1] ), .ip2(n17347), .s(n17447), .op(n16988) );
  mux2_1 U17742 ( .ip1(\x[100][0] ), .ip2(n17348), .s(n17447), .op(n16987) );
  nor2_1 U17743 ( .ip1(n17401), .ip2(n17332), .op(n17450) );
  mux2_1 U17744 ( .ip1(\x[99][15] ), .ip2(n17333), .s(n17450), .op(n16986) );
  mux2_1 U17745 ( .ip1(\x[99][14] ), .ip2(n17334), .s(n17450), .op(n16985) );
  mux2_1 U17746 ( .ip1(\x[99][13] ), .ip2(n17335), .s(n17450), .op(n16984) );
  mux2_1 U17747 ( .ip1(\x[99][12] ), .ip2(n17336), .s(n17450), .op(n16983) );
  mux2_1 U17748 ( .ip1(\x[99][11] ), .ip2(n17337), .s(n17450), .op(n16982) );
  mux2_1 U17749 ( .ip1(\x[99][10] ), .ip2(n17338), .s(n17450), .op(n16981) );
  buf_1 U17750 ( .ip(n17450), .op(n17449) );
  mux2_1 U17751 ( .ip1(\x[99][9] ), .ip2(n17339), .s(n17449), .op(n16980) );
  mux2_1 U17752 ( .ip1(\x[99][8] ), .ip2(n17340), .s(n17450), .op(n16979) );
  mux2_1 U17753 ( .ip1(\x[99][7] ), .ip2(n17341), .s(n17449), .op(n16978) );
  mux2_1 U17754 ( .ip1(\x[99][6] ), .ip2(n17342), .s(n17450), .op(n16977) );
  mux2_1 U17755 ( .ip1(\x[99][5] ), .ip2(n17343), .s(n17449), .op(n16976) );
  mux2_1 U17756 ( .ip1(\x[99][4] ), .ip2(n17344), .s(n17450), .op(n16975) );
  mux2_1 U17757 ( .ip1(\x[99][3] ), .ip2(n17345), .s(n17449), .op(n16974) );
  mux2_1 U17758 ( .ip1(\x[99][2] ), .ip2(n17346), .s(n17449), .op(n16973) );
  mux2_1 U17759 ( .ip1(\x[99][1] ), .ip2(n17347), .s(n17449), .op(n16972) );
  mux2_1 U17760 ( .ip1(\x[99][0] ), .ip2(n17348), .s(n17449), .op(n16971) );
  nor2_1 U17761 ( .ip1(n17402), .ip2(n17332), .op(n17467) );
  mux2_1 U17762 ( .ip1(\x[98][15] ), .ip2(n17333), .s(n17467), .op(n16970) );
  mux2_1 U17763 ( .ip1(\x[98][14] ), .ip2(n17334), .s(n17467), .op(n16969) );
  mux2_1 U17764 ( .ip1(\x[98][13] ), .ip2(n17335), .s(n17467), .op(n16968) );
  mux2_1 U17765 ( .ip1(\x[98][12] ), .ip2(n17336), .s(n17467), .op(n16967) );
  mux2_1 U17766 ( .ip1(\x[98][11] ), .ip2(n17337), .s(n17467), .op(n16966) );
  mux2_1 U17767 ( .ip1(\x[98][10] ), .ip2(n17338), .s(n17467), .op(n16965) );
  buf_1 U17768 ( .ip(n17467), .op(n17460) );
  mux2_1 U17769 ( .ip1(\x[98][9] ), .ip2(n17339), .s(n17460), .op(n16964) );
  mux2_1 U17770 ( .ip1(\x[98][8] ), .ip2(n17340), .s(n17467), .op(n16963) );
  mux2_1 U17771 ( .ip1(\x[98][7] ), .ip2(n17341), .s(n17460), .op(n16962) );
  mux2_1 U17772 ( .ip1(\x[98][6] ), .ip2(n17342), .s(n17467), .op(n16961) );
  mux2_1 U17773 ( .ip1(\x[98][5] ), .ip2(n17343), .s(n17460), .op(n16960) );
  mux2_1 U17774 ( .ip1(\x[98][4] ), .ip2(n17344), .s(n17467), .op(n16959) );
  mux2_1 U17775 ( .ip1(\x[98][3] ), .ip2(n17345), .s(n17460), .op(n16958) );
  mux2_1 U17776 ( .ip1(\x[98][2] ), .ip2(n17346), .s(n17460), .op(n16957) );
  mux2_1 U17777 ( .ip1(\x[98][1] ), .ip2(n17347), .s(n17460), .op(n16956) );
  mux2_1 U17778 ( .ip1(\x[98][0] ), .ip2(n17348), .s(n17460), .op(n16955) );
  nor2_1 U17779 ( .ip1(n17403), .ip2(n17332), .op(n17470) );
  mux2_1 U17780 ( .ip1(\x[97][15] ), .ip2(n17333), .s(n17470), .op(n16954) );
  mux2_1 U17781 ( .ip1(\x[97][14] ), .ip2(n17334), .s(n17470), .op(n16953) );
  mux2_1 U17782 ( .ip1(\x[97][13] ), .ip2(n17335), .s(n17470), .op(n16952) );
  mux2_1 U17783 ( .ip1(\x[97][12] ), .ip2(n17336), .s(n17470), .op(n16951) );
  mux2_1 U17784 ( .ip1(\x[97][11] ), .ip2(n17337), .s(n17470), .op(n16950) );
  mux2_1 U17785 ( .ip1(\x[97][10] ), .ip2(n17338), .s(n17470), .op(n16949) );
  buf_1 U17786 ( .ip(n17470), .op(n17469) );
  mux2_1 U17787 ( .ip1(\x[97][9] ), .ip2(n17339), .s(n17469), .op(n16948) );
  mux2_1 U17788 ( .ip1(\x[97][8] ), .ip2(n17340), .s(n17470), .op(n16947) );
  mux2_1 U17789 ( .ip1(\x[97][7] ), .ip2(n17341), .s(n17469), .op(n16946) );
  mux2_1 U17790 ( .ip1(\x[97][6] ), .ip2(n17342), .s(n17470), .op(n16945) );
  mux2_1 U17791 ( .ip1(\x[97][5] ), .ip2(n17343), .s(n17469), .op(n16944) );
  mux2_1 U17792 ( .ip1(\x[97][4] ), .ip2(n17344), .s(n17470), .op(n16943) );
  mux2_1 U17793 ( .ip1(\x[97][3] ), .ip2(n17345), .s(n17469), .op(n16942) );
  mux2_1 U17794 ( .ip1(\x[97][2] ), .ip2(n17346), .s(n17469), .op(n16941) );
  mux2_1 U17795 ( .ip1(\x[97][1] ), .ip2(n17347), .s(n17469), .op(n16940) );
  mux2_1 U17796 ( .ip1(\x[97][0] ), .ip2(n17348), .s(n17469), .op(n16939) );
  nor2_1 U17797 ( .ip1(n17405), .ip2(n17332), .op(n17472) );
  mux2_1 U17798 ( .ip1(\x[96][15] ), .ip2(n17333), .s(n17472), .op(n16938) );
  mux2_1 U17799 ( .ip1(\x[96][14] ), .ip2(n17334), .s(n17472), .op(n16937) );
  mux2_1 U17800 ( .ip1(\x[96][13] ), .ip2(n17335), .s(n17472), .op(n16936) );
  mux2_1 U17801 ( .ip1(\x[96][12] ), .ip2(n17336), .s(n17472), .op(n16935) );
  mux2_1 U17802 ( .ip1(\x[96][11] ), .ip2(n17337), .s(n17472), .op(n16934) );
  mux2_1 U17803 ( .ip1(\x[96][10] ), .ip2(n17338), .s(n17472), .op(n16933) );
  buf_1 U17804 ( .ip(n17472), .op(n17471) );
  mux2_1 U17805 ( .ip1(\x[96][9] ), .ip2(n17339), .s(n17471), .op(n16932) );
  mux2_1 U17806 ( .ip1(\x[96][8] ), .ip2(n17340), .s(n17472), .op(n16931) );
  mux2_1 U17807 ( .ip1(\x[96][7] ), .ip2(n17341), .s(n17471), .op(n16930) );
  mux2_1 U17808 ( .ip1(\x[96][6] ), .ip2(n17342), .s(n17472), .op(n16929) );
  mux2_1 U17809 ( .ip1(\x[96][5] ), .ip2(n17343), .s(n17471), .op(n16928) );
  mux2_1 U17810 ( .ip1(\x[96][4] ), .ip2(n17344), .s(n17472), .op(n16927) );
  mux2_1 U17811 ( .ip1(\x[96][3] ), .ip2(n17345), .s(n17471), .op(n16926) );
  mux2_1 U17812 ( .ip1(\x[96][2] ), .ip2(n17346), .s(n17471), .op(n16925) );
  mux2_1 U17813 ( .ip1(\x[96][1] ), .ip2(n17347), .s(n17471), .op(n16924) );
  mux2_1 U17814 ( .ip1(\x[96][0] ), .ip2(n17348), .s(n17471), .op(n16923) );
  inv_1 U17815 ( .ip(address[5]), .op(n17370) );
  nand4_1 U17816 ( .ip1(address[4]), .ip2(we), .ip3(address[6]), .ip4(n17370), 
        .op(n17349) );
  nor2_1 U17817 ( .ip1(n17373), .ip2(n17349), .op(n17474) );
  mux2_1 U17818 ( .ip1(\x[95][15] ), .ip2(n17333), .s(n17474), .op(n16922) );
  mux2_1 U17819 ( .ip1(\x[95][14] ), .ip2(n17334), .s(n17474), .op(n16921) );
  mux2_1 U17820 ( .ip1(\x[95][13] ), .ip2(n17335), .s(n17474), .op(n16920) );
  mux2_1 U17821 ( .ip1(\x[95][12] ), .ip2(n17336), .s(n17474), .op(n16919) );
  mux2_1 U17822 ( .ip1(\x[95][11] ), .ip2(n17337), .s(n17474), .op(n16918) );
  mux2_1 U17823 ( .ip1(\x[95][10] ), .ip2(n17338), .s(n17474), .op(n16917) );
  buf_1 U17824 ( .ip(n17474), .op(n17473) );
  mux2_1 U17825 ( .ip1(\x[95][9] ), .ip2(n17339), .s(n17473), .op(n16916) );
  mux2_1 U17826 ( .ip1(\x[95][8] ), .ip2(n17340), .s(n17474), .op(n16915) );
  mux2_1 U17827 ( .ip1(\x[95][7] ), .ip2(n17341), .s(n17473), .op(n16914) );
  mux2_1 U17828 ( .ip1(\x[95][6] ), .ip2(n17342), .s(n17474), .op(n16913) );
  mux2_1 U17829 ( .ip1(\x[95][5] ), .ip2(n17343), .s(n17473), .op(n16912) );
  mux2_1 U17830 ( .ip1(\x[95][4] ), .ip2(n17344), .s(n17474), .op(n16911) );
  mux2_1 U17831 ( .ip1(\x[95][3] ), .ip2(n17345), .s(n17473), .op(n16910) );
  mux2_1 U17832 ( .ip1(\x[95][2] ), .ip2(n17346), .s(n17473), .op(n16909) );
  mux2_1 U17833 ( .ip1(\x[95][1] ), .ip2(n17347), .s(n17473), .op(n16908) );
  mux2_1 U17834 ( .ip1(\x[95][0] ), .ip2(n17348), .s(n17473), .op(n16907) );
  nor2_1 U17835 ( .ip1(n17374), .ip2(n17349), .op(n17476) );
  mux2_1 U17836 ( .ip1(\x[94][15] ), .ip2(n17333), .s(n17476), .op(n16906) );
  mux2_1 U17837 ( .ip1(\x[94][14] ), .ip2(n17334), .s(n17476), .op(n16905) );
  mux2_1 U17838 ( .ip1(\x[94][13] ), .ip2(n17335), .s(n17476), .op(n16904) );
  mux2_1 U17839 ( .ip1(\x[94][12] ), .ip2(n17336), .s(n17476), .op(n16903) );
  mux2_1 U17840 ( .ip1(\x[94][11] ), .ip2(n17337), .s(n17476), .op(n16902) );
  mux2_1 U17841 ( .ip1(\x[94][10] ), .ip2(n17338), .s(n17476), .op(n16901) );
  buf_1 U17842 ( .ip(n17476), .op(n17475) );
  mux2_1 U17843 ( .ip1(\x[94][9] ), .ip2(n17339), .s(n17475), .op(n16900) );
  mux2_1 U17844 ( .ip1(\x[94][8] ), .ip2(n17340), .s(n17476), .op(n16899) );
  mux2_1 U17845 ( .ip1(\x[94][7] ), .ip2(n17341), .s(n17475), .op(n16898) );
  mux2_1 U17846 ( .ip1(\x[94][6] ), .ip2(n17342), .s(n17476), .op(n16897) );
  mux2_1 U17847 ( .ip1(\x[94][5] ), .ip2(n17343), .s(n17475), .op(n16896) );
  mux2_1 U17848 ( .ip1(\x[94][4] ), .ip2(n17344), .s(n17476), .op(n16895) );
  mux2_1 U17849 ( .ip1(\x[94][3] ), .ip2(n17345), .s(n17475), .op(n16894) );
  mux2_1 U17850 ( .ip1(\x[94][2] ), .ip2(n17346), .s(n17475), .op(n16893) );
  mux2_1 U17851 ( .ip1(\x[94][1] ), .ip2(n17347), .s(n17475), .op(n16892) );
  mux2_1 U17852 ( .ip1(\x[94][0] ), .ip2(n17348), .s(n17475), .op(n16891) );
  nor2_1 U17853 ( .ip1(n17375), .ip2(n17349), .op(n17478) );
  mux2_1 U17854 ( .ip1(\x[93][15] ), .ip2(n17333), .s(n17478), .op(n16890) );
  mux2_1 U17855 ( .ip1(\x[93][14] ), .ip2(n17334), .s(n17478), .op(n16889) );
  mux2_1 U17856 ( .ip1(\x[93][13] ), .ip2(n17335), .s(n17478), .op(n16888) );
  mux2_1 U17857 ( .ip1(\x[93][12] ), .ip2(n17336), .s(n17478), .op(n16887) );
  mux2_1 U17858 ( .ip1(\x[93][11] ), .ip2(n17337), .s(n17478), .op(n16886) );
  mux2_1 U17859 ( .ip1(\x[93][10] ), .ip2(n17338), .s(n17478), .op(n16885) );
  buf_1 U17860 ( .ip(n17478), .op(n17477) );
  mux2_1 U17861 ( .ip1(\x[93][9] ), .ip2(n17339), .s(n17477), .op(n16884) );
  mux2_1 U17862 ( .ip1(\x[93][8] ), .ip2(n17340), .s(n17478), .op(n16883) );
  mux2_1 U17863 ( .ip1(\x[93][7] ), .ip2(n17341), .s(n17477), .op(n16882) );
  mux2_1 U17864 ( .ip1(\x[93][6] ), .ip2(n17342), .s(n17478), .op(n16881) );
  mux2_1 U17865 ( .ip1(\x[93][5] ), .ip2(n17343), .s(n17477), .op(n16880) );
  mux2_1 U17866 ( .ip1(\x[93][4] ), .ip2(n17344), .s(n17478), .op(n16879) );
  mux2_1 U17867 ( .ip1(\x[93][3] ), .ip2(n17345), .s(n17477), .op(n16878) );
  mux2_1 U17868 ( .ip1(\x[93][2] ), .ip2(n17346), .s(n17477), .op(n16877) );
  mux2_1 U17869 ( .ip1(\x[93][1] ), .ip2(n17347), .s(n17477), .op(n16876) );
  mux2_1 U17870 ( .ip1(\x[93][0] ), .ip2(n17348), .s(n17477), .op(n16875) );
  nor2_1 U17871 ( .ip1(n17392), .ip2(n17349), .op(n17480) );
  mux2_1 U17872 ( .ip1(\x[92][15] ), .ip2(n17333), .s(n17480), .op(n16874) );
  mux2_1 U17873 ( .ip1(\x[92][14] ), .ip2(n17334), .s(n17480), .op(n16873) );
  mux2_1 U17874 ( .ip1(\x[92][13] ), .ip2(n17335), .s(n17480), .op(n16872) );
  mux2_1 U17875 ( .ip1(\x[92][12] ), .ip2(n17336), .s(n17480), .op(n16871) );
  mux2_1 U17876 ( .ip1(\x[92][11] ), .ip2(n17337), .s(n17480), .op(n16870) );
  mux2_1 U17877 ( .ip1(\x[92][10] ), .ip2(n17338), .s(n17480), .op(n16869) );
  buf_1 U17878 ( .ip(n17480), .op(n17479) );
  mux2_1 U17879 ( .ip1(\x[92][9] ), .ip2(n17339), .s(n17479), .op(n16868) );
  mux2_1 U17880 ( .ip1(\x[92][8] ), .ip2(n17340), .s(n17480), .op(n16867) );
  mux2_1 U17881 ( .ip1(\x[92][7] ), .ip2(n17341), .s(n17479), .op(n16866) );
  mux2_1 U17882 ( .ip1(\x[92][6] ), .ip2(n17342), .s(n17480), .op(n16865) );
  mux2_1 U17883 ( .ip1(\x[92][5] ), .ip2(n17343), .s(n17479), .op(n16864) );
  mux2_1 U17884 ( .ip1(\x[92][4] ), .ip2(n17344), .s(n17480), .op(n16863) );
  mux2_1 U17885 ( .ip1(\x[92][3] ), .ip2(n17345), .s(n17479), .op(n16862) );
  mux2_1 U17886 ( .ip1(\x[92][2] ), .ip2(n17346), .s(n17479), .op(n16861) );
  mux2_1 U17887 ( .ip1(\x[92][1] ), .ip2(n17347), .s(n17479), .op(n16860) );
  mux2_1 U17888 ( .ip1(\x[92][0] ), .ip2(n17348), .s(n17479), .op(n16859) );
  nor2_1 U17889 ( .ip1(n17393), .ip2(n17349), .op(n17482) );
  mux2_1 U17890 ( .ip1(\x[91][15] ), .ip2(n17333), .s(n17482), .op(n16858) );
  mux2_1 U17891 ( .ip1(\x[91][14] ), .ip2(n17334), .s(n17482), .op(n16857) );
  mux2_1 U17892 ( .ip1(\x[91][13] ), .ip2(n17335), .s(n17482), .op(n16856) );
  mux2_1 U17893 ( .ip1(\x[91][12] ), .ip2(n17336), .s(n17482), .op(n16855) );
  mux2_1 U17894 ( .ip1(\x[91][11] ), .ip2(n17337), .s(n17482), .op(n16854) );
  mux2_1 U17895 ( .ip1(\x[91][10] ), .ip2(n17338), .s(n17482), .op(n16853) );
  buf_1 U17896 ( .ip(n17482), .op(n17481) );
  mux2_1 U17897 ( .ip1(\x[91][9] ), .ip2(n17339), .s(n17481), .op(n16852) );
  mux2_1 U17898 ( .ip1(\x[91][8] ), .ip2(n17340), .s(n17482), .op(n16851) );
  mux2_1 U17899 ( .ip1(\x[91][7] ), .ip2(n17341), .s(n17481), .op(n16850) );
  mux2_1 U17900 ( .ip1(\x[91][6] ), .ip2(n17342), .s(n17482), .op(n16849) );
  mux2_1 U17901 ( .ip1(\x[91][5] ), .ip2(n17343), .s(n17481), .op(n16848) );
  mux2_1 U17902 ( .ip1(\x[91][4] ), .ip2(n17344), .s(n17482), .op(n16847) );
  mux2_1 U17903 ( .ip1(\x[91][3] ), .ip2(n17345), .s(n17481), .op(n16846) );
  mux2_1 U17904 ( .ip1(\x[91][2] ), .ip2(n17346), .s(n17481), .op(n16845) );
  mux2_1 U17905 ( .ip1(\x[91][1] ), .ip2(n17347), .s(n17481), .op(n16844) );
  mux2_1 U17906 ( .ip1(\x[91][0] ), .ip2(n17348), .s(n17481), .op(n16843) );
  nor2_1 U17907 ( .ip1(n17394), .ip2(n17349), .op(n17484) );
  mux2_1 U17908 ( .ip1(\x[90][15] ), .ip2(n17333), .s(n17484), .op(n16842) );
  mux2_1 U17909 ( .ip1(\x[90][14] ), .ip2(n17334), .s(n17484), .op(n16841) );
  mux2_1 U17910 ( .ip1(\x[90][13] ), .ip2(n17335), .s(n17484), .op(n16840) );
  mux2_1 U17911 ( .ip1(\x[90][12] ), .ip2(n17336), .s(n17484), .op(n16839) );
  mux2_1 U17912 ( .ip1(\x[90][11] ), .ip2(n17337), .s(n17484), .op(n16838) );
  mux2_1 U17913 ( .ip1(\x[90][10] ), .ip2(n17338), .s(n17484), .op(n16837) );
  buf_1 U17914 ( .ip(n17484), .op(n17483) );
  mux2_1 U17915 ( .ip1(\x[90][9] ), .ip2(n17339), .s(n17483), .op(n16836) );
  mux2_1 U17916 ( .ip1(\x[90][8] ), .ip2(n17340), .s(n17484), .op(n16835) );
  mux2_1 U17917 ( .ip1(\x[90][7] ), .ip2(n17341), .s(n17483), .op(n16834) );
  mux2_1 U17918 ( .ip1(\x[90][6] ), .ip2(n17342), .s(n17484), .op(n16833) );
  mux2_1 U17919 ( .ip1(\x[90][5] ), .ip2(n17343), .s(n17483), .op(n16832) );
  mux2_1 U17920 ( .ip1(\x[90][4] ), .ip2(n17344), .s(n17484), .op(n16831) );
  mux2_1 U17921 ( .ip1(\x[90][3] ), .ip2(n17345), .s(n17483), .op(n16830) );
  mux2_1 U17922 ( .ip1(\x[90][2] ), .ip2(n17346), .s(n17483), .op(n16829) );
  mux2_1 U17923 ( .ip1(\x[90][1] ), .ip2(n17347), .s(n17483), .op(n16828) );
  mux2_1 U17924 ( .ip1(\x[90][0] ), .ip2(n17348), .s(n17483), .op(n16827) );
  nor2_1 U17925 ( .ip1(n17395), .ip2(n17349), .op(n17486) );
  mux2_1 U17926 ( .ip1(\x[89][15] ), .ip2(n17333), .s(n17486), .op(n16826) );
  mux2_1 U17927 ( .ip1(\x[89][14] ), .ip2(n17334), .s(n17486), .op(n16825) );
  mux2_1 U17928 ( .ip1(\x[89][13] ), .ip2(n17335), .s(n17486), .op(n16824) );
  mux2_1 U17929 ( .ip1(\x[89][12] ), .ip2(n17336), .s(n17486), .op(n16823) );
  mux2_1 U17930 ( .ip1(\x[89][11] ), .ip2(n17337), .s(n17486), .op(n16822) );
  mux2_1 U17931 ( .ip1(\x[89][10] ), .ip2(n17338), .s(n17486), .op(n16821) );
  buf_1 U17932 ( .ip(n17486), .op(n17485) );
  mux2_1 U17933 ( .ip1(\x[89][9] ), .ip2(n17339), .s(n17485), .op(n16820) );
  mux2_1 U17934 ( .ip1(\x[89][8] ), .ip2(n17340), .s(n17486), .op(n16819) );
  mux2_1 U17935 ( .ip1(\x[89][7] ), .ip2(n17341), .s(n17485), .op(n16818) );
  mux2_1 U17936 ( .ip1(\x[89][6] ), .ip2(n17342), .s(n17486), .op(n16817) );
  mux2_1 U17937 ( .ip1(\x[89][5] ), .ip2(n17343), .s(n17485), .op(n16816) );
  mux2_1 U17938 ( .ip1(\x[89][4] ), .ip2(n17344), .s(n17486), .op(n16815) );
  mux2_1 U17939 ( .ip1(\x[89][3] ), .ip2(n17345), .s(n17485), .op(n16814) );
  mux2_1 U17940 ( .ip1(\x[89][2] ), .ip2(n17346), .s(n17485), .op(n16813) );
  mux2_1 U17941 ( .ip1(\x[89][1] ), .ip2(n17347), .s(n17485), .op(n16812) );
  mux2_1 U17942 ( .ip1(\x[89][0] ), .ip2(n17348), .s(n17485), .op(n16811) );
  nor2_1 U17943 ( .ip1(n17396), .ip2(n17349), .op(n17488) );
  mux2_1 U17944 ( .ip1(\x[88][15] ), .ip2(n17333), .s(n17488), .op(n16810) );
  mux2_1 U17945 ( .ip1(\x[88][14] ), .ip2(n17334), .s(n17488), .op(n16809) );
  mux2_1 U17946 ( .ip1(\x[88][13] ), .ip2(n17335), .s(n17488), .op(n16808) );
  mux2_1 U17947 ( .ip1(\x[88][12] ), .ip2(n17336), .s(n17488), .op(n16807) );
  mux2_1 U17948 ( .ip1(\x[88][11] ), .ip2(n17337), .s(n17488), .op(n16806) );
  mux2_1 U17949 ( .ip1(\x[88][10] ), .ip2(n17338), .s(n17488), .op(n16805) );
  buf_1 U17950 ( .ip(n17488), .op(n17487) );
  mux2_1 U17951 ( .ip1(\x[88][9] ), .ip2(n17339), .s(n17487), .op(n16804) );
  mux2_1 U17952 ( .ip1(\x[88][8] ), .ip2(n17340), .s(n17488), .op(n16803) );
  mux2_1 U17953 ( .ip1(\x[88][7] ), .ip2(n17341), .s(n17487), .op(n16802) );
  mux2_1 U17954 ( .ip1(\x[88][6] ), .ip2(n17342), .s(n17488), .op(n16801) );
  mux2_1 U17955 ( .ip1(\x[88][5] ), .ip2(n17343), .s(n17487), .op(n16800) );
  mux2_1 U17956 ( .ip1(\x[88][4] ), .ip2(n17344), .s(n17488), .op(n16799) );
  mux2_1 U17957 ( .ip1(\x[88][3] ), .ip2(n17345), .s(n17487), .op(n16798) );
  mux2_1 U17958 ( .ip1(\x[88][2] ), .ip2(n17346), .s(n17487), .op(n16797) );
  mux2_1 U17959 ( .ip1(\x[88][1] ), .ip2(n17347), .s(n17487), .op(n16796) );
  mux2_1 U17960 ( .ip1(\x[88][0] ), .ip2(n17348), .s(n17487), .op(n16795) );
  nor2_1 U17961 ( .ip1(n17397), .ip2(n17349), .op(n17490) );
  mux2_1 U17962 ( .ip1(\x[87][15] ), .ip2(n17333), .s(n17490), .op(n16794) );
  mux2_1 U17963 ( .ip1(\x[87][14] ), .ip2(n17334), .s(n17490), .op(n16793) );
  mux2_1 U17964 ( .ip1(\x[87][13] ), .ip2(n17335), .s(n17490), .op(n16792) );
  mux2_1 U17965 ( .ip1(\x[87][12] ), .ip2(n17336), .s(n17490), .op(n16791) );
  mux2_1 U17966 ( .ip1(\x[87][11] ), .ip2(n17337), .s(n17490), .op(n16790) );
  mux2_1 U17967 ( .ip1(\x[87][10] ), .ip2(n17338), .s(n17490), .op(n16789) );
  buf_1 U17968 ( .ip(n17490), .op(n17489) );
  mux2_1 U17969 ( .ip1(\x[87][9] ), .ip2(n17339), .s(n17489), .op(n16788) );
  mux2_1 U17970 ( .ip1(\x[87][8] ), .ip2(n17340), .s(n17490), .op(n16787) );
  mux2_1 U17971 ( .ip1(\x[87][7] ), .ip2(n17341), .s(n17489), .op(n16786) );
  mux2_1 U17972 ( .ip1(\x[87][6] ), .ip2(n17342), .s(n17490), .op(n16785) );
  mux2_1 U17973 ( .ip1(\x[87][5] ), .ip2(n17343), .s(n17489), .op(n16784) );
  mux2_1 U17974 ( .ip1(\x[87][4] ), .ip2(n17344), .s(n17490), .op(n16783) );
  mux2_1 U17975 ( .ip1(\x[87][3] ), .ip2(n17345), .s(n17489), .op(n16782) );
  mux2_1 U17976 ( .ip1(\x[87][2] ), .ip2(n17346), .s(n17489), .op(n16781) );
  mux2_1 U17977 ( .ip1(\x[87][1] ), .ip2(n17347), .s(n17489), .op(n16780) );
  mux2_1 U17978 ( .ip1(\x[87][0] ), .ip2(n17348), .s(n17489), .op(n16779) );
  nor2_1 U17979 ( .ip1(n17398), .ip2(n17349), .op(n17492) );
  mux2_1 U17980 ( .ip1(\x[86][15] ), .ip2(n17333), .s(n17492), .op(n16778) );
  mux2_1 U17981 ( .ip1(\x[86][14] ), .ip2(n17334), .s(n17492), .op(n16777) );
  mux2_1 U17982 ( .ip1(\x[86][13] ), .ip2(n17335), .s(n17492), .op(n16776) );
  mux2_1 U17983 ( .ip1(\x[86][12] ), .ip2(n17336), .s(n17492), .op(n16775) );
  mux2_1 U17984 ( .ip1(\x[86][11] ), .ip2(n17337), .s(n17492), .op(n16774) );
  mux2_1 U17985 ( .ip1(\x[86][10] ), .ip2(n17338), .s(n17492), .op(n16773) );
  buf_1 U17986 ( .ip(n17492), .op(n17491) );
  mux2_1 U17987 ( .ip1(\x[86][9] ), .ip2(n17339), .s(n17491), .op(n16772) );
  mux2_1 U17988 ( .ip1(\x[86][8] ), .ip2(n17340), .s(n17492), .op(n16771) );
  mux2_1 U17989 ( .ip1(\x[86][7] ), .ip2(n17341), .s(n17491), .op(n16770) );
  mux2_1 U17990 ( .ip1(\x[86][6] ), .ip2(n17342), .s(n17492), .op(n16769) );
  mux2_1 U17991 ( .ip1(\x[86][5] ), .ip2(n17343), .s(n17491), .op(n16768) );
  mux2_1 U17992 ( .ip1(\x[86][4] ), .ip2(n17344), .s(n17492), .op(n16767) );
  mux2_1 U17993 ( .ip1(\x[86][3] ), .ip2(n17345), .s(n17491), .op(n16766) );
  mux2_1 U17994 ( .ip1(\x[86][2] ), .ip2(n17346), .s(n17491), .op(n16765) );
  mux2_1 U17995 ( .ip1(\x[86][1] ), .ip2(n17347), .s(n17491), .op(n16764) );
  mux2_1 U17996 ( .ip1(\x[86][0] ), .ip2(n17348), .s(n17491), .op(n16763) );
  nor2_1 U17997 ( .ip1(n17399), .ip2(n17349), .op(n17494) );
  mux2_1 U17998 ( .ip1(\x[85][15] ), .ip2(n17333), .s(n17494), .op(n16762) );
  mux2_1 U17999 ( .ip1(\x[85][14] ), .ip2(n17334), .s(n17494), .op(n16761) );
  mux2_1 U18000 ( .ip1(\x[85][13] ), .ip2(n17335), .s(n17494), .op(n16760) );
  mux2_1 U18001 ( .ip1(\x[85][12] ), .ip2(n17336), .s(n17494), .op(n16759) );
  mux2_1 U18002 ( .ip1(\x[85][11] ), .ip2(n17337), .s(n17494), .op(n16758) );
  mux2_1 U18003 ( .ip1(\x[85][10] ), .ip2(n17338), .s(n17494), .op(n16757) );
  buf_1 U18004 ( .ip(n17494), .op(n17493) );
  mux2_1 U18005 ( .ip1(\x[85][9] ), .ip2(n17339), .s(n17493), .op(n16756) );
  mux2_1 U18006 ( .ip1(\x[85][8] ), .ip2(n17340), .s(n17494), .op(n16755) );
  mux2_1 U18007 ( .ip1(\x[85][7] ), .ip2(n17341), .s(n17493), .op(n16754) );
  mux2_1 U18008 ( .ip1(\x[85][6] ), .ip2(n17342), .s(n17494), .op(n16753) );
  mux2_1 U18009 ( .ip1(\x[85][5] ), .ip2(n17343), .s(n17493), .op(n16752) );
  mux2_1 U18010 ( .ip1(\x[85][4] ), .ip2(n17344), .s(n17494), .op(n16751) );
  mux2_1 U18011 ( .ip1(\x[85][3] ), .ip2(n17345), .s(n17493), .op(n16750) );
  mux2_1 U18012 ( .ip1(\x[85][2] ), .ip2(n17346), .s(n17493), .op(n16749) );
  mux2_1 U18013 ( .ip1(\x[85][1] ), .ip2(n17347), .s(n17493), .op(n16748) );
  mux2_1 U18014 ( .ip1(\x[85][0] ), .ip2(n17348), .s(n17493), .op(n16747) );
  buf_1 U18015 ( .ip(d[15]), .op(n17351) );
  nor2_1 U18016 ( .ip1(n17400), .ip2(n17349), .op(n17496) );
  mux2_1 U18017 ( .ip1(\x[84][15] ), .ip2(n17351), .s(n17496), .op(n16746) );
  buf_1 U18018 ( .ip(d[14]), .op(n17352) );
  mux2_1 U18019 ( .ip1(\x[84][14] ), .ip2(n17352), .s(n17496), .op(n16745) );
  buf_1 U18020 ( .ip(d[13]), .op(n17353) );
  mux2_1 U18021 ( .ip1(\x[84][13] ), .ip2(n17353), .s(n17496), .op(n16744) );
  buf_1 U18022 ( .ip(d[12]), .op(n17354) );
  mux2_1 U18023 ( .ip1(\x[84][12] ), .ip2(n17354), .s(n17496), .op(n16743) );
  buf_1 U18024 ( .ip(d[11]), .op(n17355) );
  mux2_1 U18025 ( .ip1(\x[84][11] ), .ip2(n17355), .s(n17496), .op(n16742) );
  buf_1 U18026 ( .ip(d[10]), .op(n17356) );
  mux2_1 U18027 ( .ip1(\x[84][10] ), .ip2(n17356), .s(n17496), .op(n16741) );
  buf_1 U18028 ( .ip(d[9]), .op(n17357) );
  buf_1 U18029 ( .ip(n17496), .op(n17495) );
  mux2_1 U18030 ( .ip1(\x[84][9] ), .ip2(n17357), .s(n17495), .op(n16740) );
  buf_1 U18031 ( .ip(d[8]), .op(n17358) );
  mux2_1 U18032 ( .ip1(\x[84][8] ), .ip2(n17358), .s(n17496), .op(n16739) );
  buf_1 U18033 ( .ip(d[7]), .op(n17359) );
  mux2_1 U18034 ( .ip1(\x[84][7] ), .ip2(n17359), .s(n17495), .op(n16738) );
  buf_1 U18035 ( .ip(d[6]), .op(n17360) );
  mux2_1 U18036 ( .ip1(\x[84][6] ), .ip2(n17360), .s(n17496), .op(n16737) );
  buf_1 U18037 ( .ip(d[5]), .op(n17361) );
  mux2_1 U18038 ( .ip1(\x[84][5] ), .ip2(n17361), .s(n17495), .op(n16736) );
  buf_1 U18039 ( .ip(d[4]), .op(n17362) );
  mux2_1 U18040 ( .ip1(\x[84][4] ), .ip2(n17362), .s(n17496), .op(n16735) );
  buf_1 U18041 ( .ip(d[3]), .op(n17363) );
  mux2_1 U18042 ( .ip1(\x[84][3] ), .ip2(n17363), .s(n17495), .op(n16734) );
  buf_1 U18043 ( .ip(d[2]), .op(n17364) );
  mux2_1 U18044 ( .ip1(\x[84][2] ), .ip2(n17364), .s(n17495), .op(n16733) );
  buf_1 U18045 ( .ip(d[1]), .op(n17365) );
  mux2_1 U18046 ( .ip1(\x[84][1] ), .ip2(n17365), .s(n17495), .op(n16732) );
  buf_1 U18047 ( .ip(d[0]), .op(n17366) );
  mux2_1 U18048 ( .ip1(\x[84][0] ), .ip2(n17366), .s(n17495), .op(n16731) );
  nor2_1 U18049 ( .ip1(n17401), .ip2(n17349), .op(n17498) );
  mux2_1 U18050 ( .ip1(\x[83][15] ), .ip2(n17351), .s(n17498), .op(n16730) );
  mux2_1 U18051 ( .ip1(\x[83][14] ), .ip2(n17352), .s(n17498), .op(n16729) );
  mux2_1 U18052 ( .ip1(\x[83][13] ), .ip2(n17353), .s(n17498), .op(n16728) );
  mux2_1 U18053 ( .ip1(\x[83][12] ), .ip2(n17354), .s(n17498), .op(n16727) );
  mux2_1 U18054 ( .ip1(\x[83][11] ), .ip2(n17355), .s(n17498), .op(n16726) );
  mux2_1 U18055 ( .ip1(\x[83][10] ), .ip2(n17356), .s(n17498), .op(n16725) );
  buf_1 U18056 ( .ip(n17498), .op(n17497) );
  mux2_1 U18057 ( .ip1(\x[83][9] ), .ip2(n17357), .s(n17497), .op(n16724) );
  mux2_1 U18058 ( .ip1(\x[83][8] ), .ip2(n17358), .s(n17498), .op(n16723) );
  mux2_1 U18059 ( .ip1(\x[83][7] ), .ip2(n17359), .s(n17497), .op(n16722) );
  mux2_1 U18060 ( .ip1(\x[83][6] ), .ip2(n17360), .s(n17498), .op(n16721) );
  mux2_1 U18061 ( .ip1(\x[83][5] ), .ip2(n17361), .s(n17497), .op(n16720) );
  mux2_1 U18062 ( .ip1(\x[83][4] ), .ip2(n17362), .s(n17498), .op(n16719) );
  mux2_1 U18063 ( .ip1(\x[83][3] ), .ip2(n17363), .s(n17497), .op(n16718) );
  mux2_1 U18064 ( .ip1(\x[83][2] ), .ip2(n17364), .s(n17497), .op(n16717) );
  mux2_1 U18065 ( .ip1(\x[83][1] ), .ip2(n17365), .s(n17497), .op(n16716) );
  mux2_1 U18066 ( .ip1(\x[83][0] ), .ip2(n17366), .s(n17497), .op(n16715) );
  nor2_1 U18067 ( .ip1(n17402), .ip2(n17349), .op(n17500) );
  mux2_1 U18068 ( .ip1(\x[82][15] ), .ip2(n17351), .s(n17500), .op(n16714) );
  mux2_1 U18069 ( .ip1(\x[82][14] ), .ip2(n17352), .s(n17500), .op(n16713) );
  mux2_1 U18070 ( .ip1(\x[82][13] ), .ip2(n17353), .s(n17500), .op(n16712) );
  mux2_1 U18071 ( .ip1(\x[82][12] ), .ip2(n17354), .s(n17500), .op(n16711) );
  mux2_1 U18072 ( .ip1(\x[82][11] ), .ip2(n17355), .s(n17500), .op(n16710) );
  mux2_1 U18073 ( .ip1(\x[82][10] ), .ip2(n17356), .s(n17500), .op(n16709) );
  buf_1 U18074 ( .ip(n17500), .op(n17499) );
  mux2_1 U18075 ( .ip1(\x[82][9] ), .ip2(n17357), .s(n17499), .op(n16708) );
  mux2_1 U18076 ( .ip1(\x[82][8] ), .ip2(n17358), .s(n17500), .op(n16707) );
  mux2_1 U18077 ( .ip1(\x[82][7] ), .ip2(n17359), .s(n17499), .op(n16706) );
  mux2_1 U18078 ( .ip1(\x[82][6] ), .ip2(n17360), .s(n17500), .op(n16705) );
  mux2_1 U18079 ( .ip1(\x[82][5] ), .ip2(n17361), .s(n17499), .op(n16704) );
  mux2_1 U18080 ( .ip1(\x[82][4] ), .ip2(n17362), .s(n17500), .op(n16703) );
  mux2_1 U18081 ( .ip1(\x[82][3] ), .ip2(n17363), .s(n17499), .op(n16702) );
  mux2_1 U18082 ( .ip1(\x[82][2] ), .ip2(n17364), .s(n17499), .op(n16701) );
  mux2_1 U18083 ( .ip1(\x[82][1] ), .ip2(n17365), .s(n17499), .op(n16700) );
  mux2_1 U18084 ( .ip1(\x[82][0] ), .ip2(n17366), .s(n17499), .op(n16699) );
  nor2_1 U18085 ( .ip1(n17403), .ip2(n17349), .op(n17502) );
  mux2_1 U18086 ( .ip1(\x[81][15] ), .ip2(n17351), .s(n17502), .op(n16698) );
  mux2_1 U18087 ( .ip1(\x[81][14] ), .ip2(n17352), .s(n17502), .op(n16697) );
  mux2_1 U18088 ( .ip1(\x[81][13] ), .ip2(n17353), .s(n17502), .op(n16696) );
  mux2_1 U18089 ( .ip1(\x[81][12] ), .ip2(n17354), .s(n17502), .op(n16695) );
  mux2_1 U18090 ( .ip1(\x[81][11] ), .ip2(n17355), .s(n17502), .op(n16694) );
  mux2_1 U18091 ( .ip1(\x[81][10] ), .ip2(n17356), .s(n17502), .op(n16693) );
  buf_1 U18092 ( .ip(n17502), .op(n17501) );
  mux2_1 U18093 ( .ip1(\x[81][9] ), .ip2(n17357), .s(n17501), .op(n16692) );
  mux2_1 U18094 ( .ip1(\x[81][8] ), .ip2(n17358), .s(n17502), .op(n16691) );
  mux2_1 U18095 ( .ip1(\x[81][7] ), .ip2(n17359), .s(n17501), .op(n16690) );
  mux2_1 U18096 ( .ip1(\x[81][6] ), .ip2(n17360), .s(n17502), .op(n16689) );
  mux2_1 U18097 ( .ip1(\x[81][5] ), .ip2(n17361), .s(n17501), .op(n16688) );
  mux2_1 U18098 ( .ip1(\x[81][4] ), .ip2(n17362), .s(n17502), .op(n16687) );
  mux2_1 U18099 ( .ip1(\x[81][3] ), .ip2(n17363), .s(n17501), .op(n16686) );
  mux2_1 U18100 ( .ip1(\x[81][2] ), .ip2(n17364), .s(n17501), .op(n16685) );
  mux2_1 U18101 ( .ip1(\x[81][1] ), .ip2(n17365), .s(n17501), .op(n16684) );
  mux2_1 U18102 ( .ip1(\x[81][0] ), .ip2(n17366), .s(n17501), .op(n16683) );
  nor2_1 U18103 ( .ip1(n17405), .ip2(n17349), .op(n17504) );
  mux2_1 U18104 ( .ip1(\x[80][15] ), .ip2(n17351), .s(n17504), .op(n16682) );
  mux2_1 U18105 ( .ip1(\x[80][14] ), .ip2(n17352), .s(n17504), .op(n16681) );
  mux2_1 U18106 ( .ip1(\x[80][13] ), .ip2(n17353), .s(n17504), .op(n16680) );
  mux2_1 U18107 ( .ip1(\x[80][12] ), .ip2(n17354), .s(n17504), .op(n16679) );
  mux2_1 U18108 ( .ip1(\x[80][11] ), .ip2(n17355), .s(n17504), .op(n16678) );
  mux2_1 U18109 ( .ip1(\x[80][10] ), .ip2(n17356), .s(n17504), .op(n16677) );
  buf_1 U18110 ( .ip(n17504), .op(n17503) );
  mux2_1 U18111 ( .ip1(\x[80][9] ), .ip2(n17357), .s(n17503), .op(n16676) );
  mux2_1 U18112 ( .ip1(\x[80][8] ), .ip2(n17358), .s(n17504), .op(n16675) );
  mux2_1 U18113 ( .ip1(\x[80][7] ), .ip2(n17359), .s(n17503), .op(n16674) );
  mux2_1 U18114 ( .ip1(\x[80][6] ), .ip2(n17360), .s(n17504), .op(n16673) );
  mux2_1 U18115 ( .ip1(\x[80][5] ), .ip2(n17361), .s(n17503), .op(n16672) );
  mux2_1 U18116 ( .ip1(\x[80][4] ), .ip2(n17362), .s(n17504), .op(n16671) );
  mux2_1 U18117 ( .ip1(\x[80][3] ), .ip2(n17363), .s(n17503), .op(n16670) );
  mux2_1 U18118 ( .ip1(\x[80][2] ), .ip2(n17364), .s(n17503), .op(n16669) );
  mux2_1 U18119 ( .ip1(\x[80][1] ), .ip2(n17365), .s(n17503), .op(n16668) );
  mux2_1 U18120 ( .ip1(\x[80][0] ), .ip2(n17366), .s(n17503), .op(n16667) );
  nand3_1 U18121 ( .ip1(address[6]), .ip2(n17372), .ip3(n17370), .op(n17350)
         );
  nor2_1 U18122 ( .ip1(n17373), .ip2(n17350), .op(n17506) );
  mux2_1 U18123 ( .ip1(\x[79][15] ), .ip2(n17351), .s(n17506), .op(n16666) );
  mux2_1 U18124 ( .ip1(\x[79][14] ), .ip2(n17352), .s(n17506), .op(n16665) );
  mux2_1 U18125 ( .ip1(\x[79][13] ), .ip2(n17353), .s(n17506), .op(n16664) );
  mux2_1 U18126 ( .ip1(\x[79][12] ), .ip2(n17354), .s(n17506), .op(n16663) );
  mux2_1 U18127 ( .ip1(\x[79][11] ), .ip2(n17355), .s(n17506), .op(n16662) );
  mux2_1 U18128 ( .ip1(\x[79][10] ), .ip2(n17356), .s(n17506), .op(n16661) );
  buf_1 U18129 ( .ip(n17506), .op(n17505) );
  mux2_1 U18130 ( .ip1(\x[79][9] ), .ip2(n17357), .s(n17505), .op(n16660) );
  mux2_1 U18131 ( .ip1(\x[79][8] ), .ip2(n17358), .s(n17506), .op(n16659) );
  mux2_1 U18132 ( .ip1(\x[79][7] ), .ip2(n17359), .s(n17505), .op(n16658) );
  mux2_1 U18133 ( .ip1(\x[79][6] ), .ip2(n17360), .s(n17506), .op(n16657) );
  mux2_1 U18134 ( .ip1(\x[79][5] ), .ip2(n17361), .s(n17505), .op(n16656) );
  mux2_1 U18135 ( .ip1(\x[79][4] ), .ip2(n17362), .s(n17506), .op(n16655) );
  mux2_1 U18136 ( .ip1(\x[79][3] ), .ip2(n17363), .s(n17505), .op(n16654) );
  mux2_1 U18137 ( .ip1(\x[79][2] ), .ip2(n17364), .s(n17505), .op(n16653) );
  mux2_1 U18138 ( .ip1(\x[79][1] ), .ip2(n17365), .s(n17505), .op(n16652) );
  mux2_1 U18139 ( .ip1(\x[79][0] ), .ip2(n17366), .s(n17505), .op(n16651) );
  nor2_1 U18140 ( .ip1(n17374), .ip2(n17350), .op(n17508) );
  mux2_1 U18141 ( .ip1(\x[78][15] ), .ip2(n17351), .s(n17508), .op(n16650) );
  mux2_1 U18142 ( .ip1(\x[78][14] ), .ip2(n17352), .s(n17508), .op(n16649) );
  mux2_1 U18143 ( .ip1(\x[78][13] ), .ip2(n17353), .s(n17508), .op(n16648) );
  mux2_1 U18144 ( .ip1(\x[78][12] ), .ip2(n17354), .s(n17508), .op(n16647) );
  mux2_1 U18145 ( .ip1(\x[78][11] ), .ip2(n17355), .s(n17508), .op(n16646) );
  mux2_1 U18146 ( .ip1(\x[78][10] ), .ip2(n17356), .s(n17508), .op(n16645) );
  buf_1 U18147 ( .ip(n17508), .op(n17507) );
  mux2_1 U18148 ( .ip1(\x[78][9] ), .ip2(n17357), .s(n17507), .op(n16644) );
  mux2_1 U18149 ( .ip1(\x[78][8] ), .ip2(n17358), .s(n17508), .op(n16643) );
  mux2_1 U18150 ( .ip1(\x[78][7] ), .ip2(n17359), .s(n17507), .op(n16642) );
  mux2_1 U18151 ( .ip1(\x[78][6] ), .ip2(n17360), .s(n17508), .op(n16641) );
  mux2_1 U18152 ( .ip1(\x[78][5] ), .ip2(n17361), .s(n17507), .op(n16640) );
  mux2_1 U18153 ( .ip1(\x[78][4] ), .ip2(n17362), .s(n17508), .op(n16639) );
  mux2_1 U18154 ( .ip1(\x[78][3] ), .ip2(n17363), .s(n17507), .op(n16638) );
  mux2_1 U18155 ( .ip1(\x[78][2] ), .ip2(n17364), .s(n17507), .op(n16637) );
  mux2_1 U18156 ( .ip1(\x[78][1] ), .ip2(n17365), .s(n17507), .op(n16636) );
  mux2_1 U18157 ( .ip1(\x[78][0] ), .ip2(n17366), .s(n17507), .op(n16635) );
  nor2_1 U18158 ( .ip1(n17375), .ip2(n17350), .op(n17510) );
  mux2_1 U18159 ( .ip1(\x[77][15] ), .ip2(n17351), .s(n17510), .op(n16634) );
  mux2_1 U18160 ( .ip1(\x[77][14] ), .ip2(n17352), .s(n17510), .op(n16633) );
  mux2_1 U18161 ( .ip1(\x[77][13] ), .ip2(n17353), .s(n17510), .op(n16632) );
  mux2_1 U18162 ( .ip1(\x[77][12] ), .ip2(n17354), .s(n17510), .op(n16631) );
  mux2_1 U18163 ( .ip1(\x[77][11] ), .ip2(n17355), .s(n17510), .op(n16630) );
  mux2_1 U18164 ( .ip1(\x[77][10] ), .ip2(n17356), .s(n17510), .op(n16629) );
  buf_1 U18165 ( .ip(n17510), .op(n17509) );
  mux2_1 U18166 ( .ip1(\x[77][9] ), .ip2(n17357), .s(n17509), .op(n16628) );
  mux2_1 U18167 ( .ip1(\x[77][8] ), .ip2(n17358), .s(n17510), .op(n16627) );
  mux2_1 U18168 ( .ip1(\x[77][7] ), .ip2(n17359), .s(n17509), .op(n16626) );
  mux2_1 U18169 ( .ip1(\x[77][6] ), .ip2(n17360), .s(n17510), .op(n16625) );
  mux2_1 U18170 ( .ip1(\x[77][5] ), .ip2(n17361), .s(n17509), .op(n16624) );
  mux2_1 U18171 ( .ip1(\x[77][4] ), .ip2(n17362), .s(n17510), .op(n16623) );
  mux2_1 U18172 ( .ip1(\x[77][3] ), .ip2(n17363), .s(n17509), .op(n16622) );
  mux2_1 U18173 ( .ip1(\x[77][2] ), .ip2(n17364), .s(n17509), .op(n16621) );
  mux2_1 U18174 ( .ip1(\x[77][1] ), .ip2(n17365), .s(n17509), .op(n16620) );
  mux2_1 U18175 ( .ip1(\x[77][0] ), .ip2(n17366), .s(n17509), .op(n16619) );
  nor2_1 U18176 ( .ip1(n17392), .ip2(n17350), .op(n17512) );
  mux2_1 U18177 ( .ip1(\x[76][15] ), .ip2(n17351), .s(n17512), .op(n16618) );
  mux2_1 U18178 ( .ip1(\x[76][14] ), .ip2(n17352), .s(n17512), .op(n16617) );
  mux2_1 U18179 ( .ip1(\x[76][13] ), .ip2(n17353), .s(n17512), .op(n16616) );
  mux2_1 U18180 ( .ip1(\x[76][12] ), .ip2(n17354), .s(n17512), .op(n16615) );
  mux2_1 U18181 ( .ip1(\x[76][11] ), .ip2(n17355), .s(n17512), .op(n16614) );
  mux2_1 U18182 ( .ip1(\x[76][10] ), .ip2(n17356), .s(n17512), .op(n16613) );
  buf_1 U18183 ( .ip(n17512), .op(n17511) );
  mux2_1 U18184 ( .ip1(\x[76][9] ), .ip2(n17357), .s(n17511), .op(n16612) );
  mux2_1 U18185 ( .ip1(\x[76][8] ), .ip2(n17358), .s(n17512), .op(n16611) );
  mux2_1 U18186 ( .ip1(\x[76][7] ), .ip2(n17359), .s(n17511), .op(n16610) );
  mux2_1 U18187 ( .ip1(\x[76][6] ), .ip2(n17360), .s(n17512), .op(n16609) );
  mux2_1 U18188 ( .ip1(\x[76][5] ), .ip2(n17361), .s(n17511), .op(n16608) );
  mux2_1 U18189 ( .ip1(\x[76][4] ), .ip2(n17362), .s(n17512), .op(n16607) );
  mux2_1 U18190 ( .ip1(\x[76][3] ), .ip2(n17363), .s(n17511), .op(n16606) );
  mux2_1 U18191 ( .ip1(\x[76][2] ), .ip2(n17364), .s(n17511), .op(n16605) );
  mux2_1 U18192 ( .ip1(\x[76][1] ), .ip2(n17365), .s(n17511), .op(n16604) );
  mux2_1 U18193 ( .ip1(\x[76][0] ), .ip2(n17366), .s(n17511), .op(n16603) );
  nor2_1 U18194 ( .ip1(n17393), .ip2(n17350), .op(n17514) );
  mux2_1 U18195 ( .ip1(\x[75][15] ), .ip2(n17351), .s(n17514), .op(n16602) );
  mux2_1 U18196 ( .ip1(\x[75][14] ), .ip2(n17352), .s(n17514), .op(n16601) );
  mux2_1 U18197 ( .ip1(\x[75][13] ), .ip2(n17353), .s(n17514), .op(n16600) );
  mux2_1 U18198 ( .ip1(\x[75][12] ), .ip2(n17354), .s(n17514), .op(n16599) );
  mux2_1 U18199 ( .ip1(\x[75][11] ), .ip2(n17355), .s(n17514), .op(n16598) );
  mux2_1 U18200 ( .ip1(\x[75][10] ), .ip2(n17356), .s(n17514), .op(n16597) );
  buf_1 U18201 ( .ip(n17514), .op(n17513) );
  mux2_1 U18202 ( .ip1(\x[75][9] ), .ip2(n17357), .s(n17513), .op(n16596) );
  mux2_1 U18203 ( .ip1(\x[75][8] ), .ip2(n17358), .s(n17514), .op(n16595) );
  mux2_1 U18204 ( .ip1(\x[75][7] ), .ip2(n17359), .s(n17513), .op(n16594) );
  mux2_1 U18205 ( .ip1(\x[75][6] ), .ip2(n17360), .s(n17514), .op(n16593) );
  mux2_1 U18206 ( .ip1(\x[75][5] ), .ip2(n17361), .s(n17513), .op(n16592) );
  mux2_1 U18207 ( .ip1(\x[75][4] ), .ip2(n17362), .s(n17514), .op(n16591) );
  mux2_1 U18208 ( .ip1(\x[75][3] ), .ip2(n17363), .s(n17513), .op(n16590) );
  mux2_1 U18209 ( .ip1(\x[75][2] ), .ip2(n17364), .s(n17513), .op(n16589) );
  mux2_1 U18210 ( .ip1(\x[75][1] ), .ip2(n17365), .s(n17513), .op(n16588) );
  mux2_1 U18211 ( .ip1(\x[75][0] ), .ip2(n17366), .s(n17513), .op(n16587) );
  nor2_1 U18212 ( .ip1(n17394), .ip2(n17350), .op(n17516) );
  mux2_1 U18213 ( .ip1(\x[74][15] ), .ip2(n17351), .s(n17516), .op(n16586) );
  mux2_1 U18214 ( .ip1(\x[74][14] ), .ip2(n17352), .s(n17516), .op(n16585) );
  mux2_1 U18215 ( .ip1(\x[74][13] ), .ip2(n17353), .s(n17516), .op(n16584) );
  mux2_1 U18216 ( .ip1(\x[74][12] ), .ip2(n17354), .s(n17516), .op(n16583) );
  mux2_1 U18217 ( .ip1(\x[74][11] ), .ip2(n17355), .s(n17516), .op(n16582) );
  mux2_1 U18218 ( .ip1(\x[74][10] ), .ip2(n17356), .s(n17516), .op(n16581) );
  buf_1 U18219 ( .ip(n17516), .op(n17515) );
  mux2_1 U18220 ( .ip1(\x[74][9] ), .ip2(n17357), .s(n17515), .op(n16580) );
  mux2_1 U18221 ( .ip1(\x[74][8] ), .ip2(n17358), .s(n17516), .op(n16579) );
  mux2_1 U18222 ( .ip1(\x[74][7] ), .ip2(n17359), .s(n17515), .op(n16578) );
  mux2_1 U18223 ( .ip1(\x[74][6] ), .ip2(n17360), .s(n17516), .op(n16577) );
  mux2_1 U18224 ( .ip1(\x[74][5] ), .ip2(n17361), .s(n17515), .op(n16576) );
  mux2_1 U18225 ( .ip1(\x[74][4] ), .ip2(n17362), .s(n17516), .op(n16575) );
  mux2_1 U18226 ( .ip1(\x[74][3] ), .ip2(n17363), .s(n17515), .op(n16574) );
  mux2_1 U18227 ( .ip1(\x[74][2] ), .ip2(n17364), .s(n17515), .op(n16573) );
  mux2_1 U18228 ( .ip1(\x[74][1] ), .ip2(n17365), .s(n17515), .op(n16572) );
  mux2_1 U18229 ( .ip1(\x[74][0] ), .ip2(n17366), .s(n17515), .op(n16571) );
  nor2_1 U18230 ( .ip1(n17395), .ip2(n17350), .op(n17518) );
  mux2_1 U18231 ( .ip1(\x[73][15] ), .ip2(n17351), .s(n17518), .op(n16570) );
  mux2_1 U18232 ( .ip1(\x[73][14] ), .ip2(n17352), .s(n17518), .op(n16569) );
  mux2_1 U18233 ( .ip1(\x[73][13] ), .ip2(n17353), .s(n17518), .op(n16568) );
  mux2_1 U18234 ( .ip1(\x[73][12] ), .ip2(n17354), .s(n17518), .op(n16567) );
  mux2_1 U18235 ( .ip1(\x[73][11] ), .ip2(n17355), .s(n17518), .op(n16566) );
  mux2_1 U18236 ( .ip1(\x[73][10] ), .ip2(n17356), .s(n17518), .op(n16565) );
  buf_1 U18237 ( .ip(n17518), .op(n17517) );
  mux2_1 U18238 ( .ip1(\x[73][9] ), .ip2(n17357), .s(n17517), .op(n16564) );
  mux2_1 U18239 ( .ip1(\x[73][8] ), .ip2(n17358), .s(n17518), .op(n16563) );
  mux2_1 U18240 ( .ip1(\x[73][7] ), .ip2(n17359), .s(n17517), .op(n16562) );
  mux2_1 U18241 ( .ip1(\x[73][6] ), .ip2(n17360), .s(n17518), .op(n16561) );
  mux2_1 U18242 ( .ip1(\x[73][5] ), .ip2(n17361), .s(n17517), .op(n16560) );
  mux2_1 U18243 ( .ip1(\x[73][4] ), .ip2(n17362), .s(n17518), .op(n16559) );
  mux2_1 U18244 ( .ip1(\x[73][3] ), .ip2(n17363), .s(n17517), .op(n16558) );
  mux2_1 U18245 ( .ip1(\x[73][2] ), .ip2(n17364), .s(n17517), .op(n16557) );
  mux2_1 U18246 ( .ip1(\x[73][1] ), .ip2(n17365), .s(n17517), .op(n16556) );
  mux2_1 U18247 ( .ip1(\x[73][0] ), .ip2(n17366), .s(n17517), .op(n16555) );
  nor2_1 U18248 ( .ip1(n17396), .ip2(n17350), .op(n17520) );
  mux2_1 U18249 ( .ip1(\x[72][15] ), .ip2(n17351), .s(n17520), .op(n16554) );
  mux2_1 U18250 ( .ip1(\x[72][14] ), .ip2(n17352), .s(n17520), .op(n16553) );
  mux2_1 U18251 ( .ip1(\x[72][13] ), .ip2(n17353), .s(n17520), .op(n16552) );
  mux2_1 U18252 ( .ip1(\x[72][12] ), .ip2(n17354), .s(n17520), .op(n16551) );
  mux2_1 U18253 ( .ip1(\x[72][11] ), .ip2(n17355), .s(n17520), .op(n16550) );
  mux2_1 U18254 ( .ip1(\x[72][10] ), .ip2(n17356), .s(n17520), .op(n16549) );
  buf_1 U18255 ( .ip(n17520), .op(n17519) );
  mux2_1 U18256 ( .ip1(\x[72][9] ), .ip2(n17357), .s(n17519), .op(n16548) );
  mux2_1 U18257 ( .ip1(\x[72][8] ), .ip2(n17358), .s(n17520), .op(n16547) );
  mux2_1 U18258 ( .ip1(\x[72][7] ), .ip2(n17359), .s(n17519), .op(n16546) );
  mux2_1 U18259 ( .ip1(\x[72][6] ), .ip2(n17360), .s(n17520), .op(n16545) );
  mux2_1 U18260 ( .ip1(\x[72][5] ), .ip2(n17361), .s(n17519), .op(n16544) );
  mux2_1 U18261 ( .ip1(\x[72][4] ), .ip2(n17362), .s(n17520), .op(n16543) );
  mux2_1 U18262 ( .ip1(\x[72][3] ), .ip2(n17363), .s(n17519), .op(n16542) );
  mux2_1 U18263 ( .ip1(\x[72][2] ), .ip2(n17364), .s(n17519), .op(n16541) );
  mux2_1 U18264 ( .ip1(\x[72][1] ), .ip2(n17365), .s(n17519), .op(n16540) );
  mux2_1 U18265 ( .ip1(\x[72][0] ), .ip2(n17366), .s(n17519), .op(n16539) );
  nor2_1 U18266 ( .ip1(n17397), .ip2(n17350), .op(n17522) );
  mux2_1 U18267 ( .ip1(\x[71][15] ), .ip2(n17351), .s(n17522), .op(n16538) );
  mux2_1 U18268 ( .ip1(\x[71][14] ), .ip2(n17352), .s(n17522), .op(n16537) );
  mux2_1 U18269 ( .ip1(\x[71][13] ), .ip2(n17353), .s(n17522), .op(n16536) );
  mux2_1 U18270 ( .ip1(\x[71][12] ), .ip2(n17354), .s(n17522), .op(n16535) );
  mux2_1 U18271 ( .ip1(\x[71][11] ), .ip2(n17355), .s(n17522), .op(n16534) );
  mux2_1 U18272 ( .ip1(\x[71][10] ), .ip2(n17356), .s(n17522), .op(n16533) );
  buf_1 U18273 ( .ip(n17522), .op(n17521) );
  mux2_1 U18274 ( .ip1(\x[71][9] ), .ip2(n17357), .s(n17521), .op(n16532) );
  mux2_1 U18275 ( .ip1(\x[71][8] ), .ip2(n17358), .s(n17522), .op(n16531) );
  mux2_1 U18276 ( .ip1(\x[71][7] ), .ip2(n17359), .s(n17521), .op(n16530) );
  mux2_1 U18277 ( .ip1(\x[71][6] ), .ip2(n17360), .s(n17522), .op(n16529) );
  mux2_1 U18278 ( .ip1(\x[71][5] ), .ip2(n17361), .s(n17521), .op(n16528) );
  mux2_1 U18279 ( .ip1(\x[71][4] ), .ip2(n17362), .s(n17522), .op(n16527) );
  mux2_1 U18280 ( .ip1(\x[71][3] ), .ip2(n17363), .s(n17521), .op(n16526) );
  mux2_1 U18281 ( .ip1(\x[71][2] ), .ip2(n17364), .s(n17521), .op(n16525) );
  mux2_1 U18282 ( .ip1(\x[71][1] ), .ip2(n17365), .s(n17521), .op(n16524) );
  mux2_1 U18283 ( .ip1(\x[71][0] ), .ip2(n17366), .s(n17521), .op(n16523) );
  nor2_1 U18284 ( .ip1(n17398), .ip2(n17350), .op(n17524) );
  mux2_1 U18285 ( .ip1(\x[70][15] ), .ip2(n17351), .s(n17524), .op(n16522) );
  mux2_1 U18286 ( .ip1(\x[70][14] ), .ip2(n17352), .s(n17524), .op(n16521) );
  mux2_1 U18287 ( .ip1(\x[70][13] ), .ip2(n17353), .s(n17524), .op(n16520) );
  mux2_1 U18288 ( .ip1(\x[70][12] ), .ip2(n17354), .s(n17524), .op(n16519) );
  mux2_1 U18289 ( .ip1(\x[70][11] ), .ip2(n17355), .s(n17524), .op(n16518) );
  mux2_1 U18290 ( .ip1(\x[70][10] ), .ip2(n17356), .s(n17524), .op(n16517) );
  buf_1 U18291 ( .ip(n17524), .op(n17523) );
  mux2_1 U18292 ( .ip1(\x[70][9] ), .ip2(n17357), .s(n17523), .op(n16516) );
  mux2_1 U18293 ( .ip1(\x[70][8] ), .ip2(n17358), .s(n17524), .op(n16515) );
  mux2_1 U18294 ( .ip1(\x[70][7] ), .ip2(n17359), .s(n17523), .op(n16514) );
  mux2_1 U18295 ( .ip1(\x[70][6] ), .ip2(n17360), .s(n17524), .op(n16513) );
  mux2_1 U18296 ( .ip1(\x[70][5] ), .ip2(n17361), .s(n17523), .op(n16512) );
  mux2_1 U18297 ( .ip1(\x[70][4] ), .ip2(n17362), .s(n17524), .op(n16511) );
  mux2_1 U18298 ( .ip1(\x[70][3] ), .ip2(n17363), .s(n17523), .op(n16510) );
  mux2_1 U18299 ( .ip1(\x[70][2] ), .ip2(n17364), .s(n17523), .op(n16509) );
  mux2_1 U18300 ( .ip1(\x[70][1] ), .ip2(n17365), .s(n17523), .op(n16508) );
  mux2_1 U18301 ( .ip1(\x[70][0] ), .ip2(n17366), .s(n17523), .op(n16507) );
  nor2_1 U18302 ( .ip1(n17399), .ip2(n17350), .op(n17526) );
  mux2_1 U18303 ( .ip1(\x[69][15] ), .ip2(n17351), .s(n17526), .op(n16506) );
  mux2_1 U18304 ( .ip1(\x[69][14] ), .ip2(n17352), .s(n17526), .op(n16505) );
  mux2_1 U18305 ( .ip1(\x[69][13] ), .ip2(n17353), .s(n17526), .op(n16504) );
  mux2_1 U18306 ( .ip1(\x[69][12] ), .ip2(n17354), .s(n17526), .op(n16503) );
  mux2_1 U18307 ( .ip1(\x[69][11] ), .ip2(n17355), .s(n17526), .op(n16502) );
  mux2_1 U18308 ( .ip1(\x[69][10] ), .ip2(n17356), .s(n17526), .op(n16501) );
  buf_1 U18309 ( .ip(n17526), .op(n17525) );
  mux2_1 U18310 ( .ip1(\x[69][9] ), .ip2(n17357), .s(n17525), .op(n16500) );
  mux2_1 U18311 ( .ip1(\x[69][8] ), .ip2(n17358), .s(n17526), .op(n16499) );
  mux2_1 U18312 ( .ip1(\x[69][7] ), .ip2(n17359), .s(n17525), .op(n16498) );
  mux2_1 U18313 ( .ip1(\x[69][6] ), .ip2(n17360), .s(n17526), .op(n16497) );
  mux2_1 U18314 ( .ip1(\x[69][5] ), .ip2(n17361), .s(n17525), .op(n16496) );
  mux2_1 U18315 ( .ip1(\x[69][4] ), .ip2(n17362), .s(n17526), .op(n16495) );
  mux2_1 U18316 ( .ip1(\x[69][3] ), .ip2(n17363), .s(n17525), .op(n16494) );
  mux2_1 U18317 ( .ip1(\x[69][2] ), .ip2(n17364), .s(n17525), .op(n16493) );
  mux2_1 U18318 ( .ip1(\x[69][1] ), .ip2(n17365), .s(n17525), .op(n16492) );
  mux2_1 U18319 ( .ip1(\x[69][0] ), .ip2(n17366), .s(n17525), .op(n16491) );
  nor2_1 U18320 ( .ip1(n17400), .ip2(n17350), .op(n17528) );
  mux2_1 U18321 ( .ip1(\x[68][15] ), .ip2(n17351), .s(n17528), .op(n16490) );
  mux2_1 U18322 ( .ip1(\x[68][14] ), .ip2(n17352), .s(n17528), .op(n16489) );
  mux2_1 U18323 ( .ip1(\x[68][13] ), .ip2(n17353), .s(n17528), .op(n16488) );
  mux2_1 U18324 ( .ip1(\x[68][12] ), .ip2(n17354), .s(n17528), .op(n16487) );
  mux2_1 U18325 ( .ip1(\x[68][11] ), .ip2(n17355), .s(n17528), .op(n16486) );
  mux2_1 U18326 ( .ip1(\x[68][10] ), .ip2(n17356), .s(n17528), .op(n16485) );
  buf_1 U18327 ( .ip(n17528), .op(n17527) );
  mux2_1 U18328 ( .ip1(\x[68][9] ), .ip2(n17357), .s(n17527), .op(n16484) );
  mux2_1 U18329 ( .ip1(\x[68][8] ), .ip2(n17358), .s(n17528), .op(n16483) );
  mux2_1 U18330 ( .ip1(\x[68][7] ), .ip2(n17359), .s(n17527), .op(n16482) );
  mux2_1 U18331 ( .ip1(\x[68][6] ), .ip2(n17360), .s(n17528), .op(n16481) );
  mux2_1 U18332 ( .ip1(\x[68][5] ), .ip2(n17361), .s(n17527), .op(n16480) );
  mux2_1 U18333 ( .ip1(\x[68][4] ), .ip2(n17362), .s(n17528), .op(n16479) );
  mux2_1 U18334 ( .ip1(\x[68][3] ), .ip2(n17363), .s(n17527), .op(n16478) );
  mux2_1 U18335 ( .ip1(\x[68][2] ), .ip2(n17364), .s(n17527), .op(n16477) );
  mux2_1 U18336 ( .ip1(\x[68][1] ), .ip2(n17365), .s(n17527), .op(n16476) );
  mux2_1 U18337 ( .ip1(\x[68][0] ), .ip2(n17366), .s(n17527), .op(n16475) );
  nor2_1 U18338 ( .ip1(n17401), .ip2(n17350), .op(n17530) );
  mux2_1 U18339 ( .ip1(\x[67][15] ), .ip2(n17351), .s(n17530), .op(n16474) );
  mux2_1 U18340 ( .ip1(\x[67][14] ), .ip2(n17352), .s(n17530), .op(n16473) );
  mux2_1 U18341 ( .ip1(\x[67][13] ), .ip2(n17353), .s(n17530), .op(n16472) );
  mux2_1 U18342 ( .ip1(\x[67][12] ), .ip2(n17354), .s(n17530), .op(n16471) );
  mux2_1 U18343 ( .ip1(\x[67][11] ), .ip2(n17355), .s(n17530), .op(n16470) );
  mux2_1 U18344 ( .ip1(\x[67][10] ), .ip2(n17356), .s(n17530), .op(n16469) );
  buf_1 U18345 ( .ip(n17530), .op(n17529) );
  mux2_1 U18346 ( .ip1(\x[67][9] ), .ip2(n17357), .s(n17529), .op(n16468) );
  mux2_1 U18347 ( .ip1(\x[67][8] ), .ip2(n17358), .s(n17530), .op(n16467) );
  mux2_1 U18348 ( .ip1(\x[67][7] ), .ip2(n17359), .s(n17529), .op(n16466) );
  mux2_1 U18349 ( .ip1(\x[67][6] ), .ip2(n17360), .s(n17530), .op(n16465) );
  mux2_1 U18350 ( .ip1(\x[67][5] ), .ip2(n17361), .s(n17529), .op(n16464) );
  mux2_1 U18351 ( .ip1(\x[67][4] ), .ip2(n17362), .s(n17530), .op(n16463) );
  mux2_1 U18352 ( .ip1(\x[67][3] ), .ip2(n17363), .s(n17529), .op(n16462) );
  mux2_1 U18353 ( .ip1(\x[67][2] ), .ip2(n17364), .s(n17529), .op(n16461) );
  mux2_1 U18354 ( .ip1(\x[67][1] ), .ip2(n17365), .s(n17529), .op(n16460) );
  mux2_1 U18355 ( .ip1(\x[67][0] ), .ip2(n17366), .s(n17529), .op(n16459) );
  nor2_1 U18356 ( .ip1(n17402), .ip2(n17350), .op(n17532) );
  mux2_1 U18357 ( .ip1(\x[66][15] ), .ip2(n17351), .s(n17532), .op(n16458) );
  mux2_1 U18358 ( .ip1(\x[66][14] ), .ip2(n17352), .s(n17532), .op(n16457) );
  mux2_1 U18359 ( .ip1(\x[66][13] ), .ip2(n17353), .s(n17532), .op(n16456) );
  mux2_1 U18360 ( .ip1(\x[66][12] ), .ip2(n17354), .s(n17532), .op(n16455) );
  mux2_1 U18361 ( .ip1(\x[66][11] ), .ip2(n17355), .s(n17532), .op(n16454) );
  mux2_1 U18362 ( .ip1(\x[66][10] ), .ip2(n17356), .s(n17532), .op(n16453) );
  buf_1 U18363 ( .ip(n17532), .op(n17531) );
  mux2_1 U18364 ( .ip1(\x[66][9] ), .ip2(n17357), .s(n17531), .op(n16452) );
  mux2_1 U18365 ( .ip1(\x[66][8] ), .ip2(n17358), .s(n17532), .op(n16451) );
  mux2_1 U18366 ( .ip1(\x[66][7] ), .ip2(n17359), .s(n17531), .op(n16450) );
  mux2_1 U18367 ( .ip1(\x[66][6] ), .ip2(n17360), .s(n17532), .op(n16449) );
  mux2_1 U18368 ( .ip1(\x[66][5] ), .ip2(n17361), .s(n17531), .op(n16448) );
  mux2_1 U18369 ( .ip1(\x[66][4] ), .ip2(n17362), .s(n17532), .op(n16447) );
  mux2_1 U18370 ( .ip1(\x[66][3] ), .ip2(n17363), .s(n17531), .op(n16446) );
  mux2_1 U18371 ( .ip1(\x[66][2] ), .ip2(n17364), .s(n17531), .op(n16445) );
  mux2_1 U18372 ( .ip1(\x[66][1] ), .ip2(n17365), .s(n17531), .op(n16444) );
  mux2_1 U18373 ( .ip1(\x[66][0] ), .ip2(n17366), .s(n17531), .op(n16443) );
  nor2_1 U18374 ( .ip1(n17403), .ip2(n17350), .op(n17534) );
  mux2_1 U18375 ( .ip1(\x[65][15] ), .ip2(n17351), .s(n17534), .op(n16442) );
  mux2_1 U18376 ( .ip1(\x[65][14] ), .ip2(n17352), .s(n17534), .op(n16441) );
  mux2_1 U18377 ( .ip1(\x[65][13] ), .ip2(n17353), .s(n17534), .op(n16440) );
  mux2_1 U18378 ( .ip1(\x[65][12] ), .ip2(n17354), .s(n17534), .op(n16439) );
  mux2_1 U18379 ( .ip1(\x[65][11] ), .ip2(n17355), .s(n17534), .op(n16438) );
  mux2_1 U18380 ( .ip1(\x[65][10] ), .ip2(n17356), .s(n17534), .op(n16437) );
  buf_1 U18381 ( .ip(n17534), .op(n17533) );
  mux2_1 U18382 ( .ip1(\x[65][9] ), .ip2(n17357), .s(n17533), .op(n16436) );
  mux2_1 U18383 ( .ip1(\x[65][8] ), .ip2(n17358), .s(n17534), .op(n16435) );
  mux2_1 U18384 ( .ip1(\x[65][7] ), .ip2(n17359), .s(n17533), .op(n16434) );
  mux2_1 U18385 ( .ip1(\x[65][6] ), .ip2(n17360), .s(n17534), .op(n16433) );
  mux2_1 U18386 ( .ip1(\x[65][5] ), .ip2(n17361), .s(n17533), .op(n16432) );
  mux2_1 U18387 ( .ip1(\x[65][4] ), .ip2(n17362), .s(n17534), .op(n16431) );
  mux2_1 U18388 ( .ip1(\x[65][3] ), .ip2(n17363), .s(n17533), .op(n16430) );
  mux2_1 U18389 ( .ip1(\x[65][2] ), .ip2(n17364), .s(n17533), .op(n16429) );
  mux2_1 U18390 ( .ip1(\x[65][1] ), .ip2(n17365), .s(n17533), .op(n16428) );
  mux2_1 U18391 ( .ip1(\x[65][0] ), .ip2(n17366), .s(n17533), .op(n16427) );
  nor2_1 U18392 ( .ip1(n17405), .ip2(n17350), .op(n17536) );
  mux2_1 U18393 ( .ip1(\x[64][15] ), .ip2(n17351), .s(n17536), .op(n16426) );
  mux2_1 U18394 ( .ip1(\x[64][14] ), .ip2(n17352), .s(n17536), .op(n16425) );
  mux2_1 U18395 ( .ip1(\x[64][13] ), .ip2(n17353), .s(n17536), .op(n16424) );
  mux2_1 U18396 ( .ip1(\x[64][12] ), .ip2(n17354), .s(n17536), .op(n16423) );
  mux2_1 U18397 ( .ip1(\x[64][11] ), .ip2(n17355), .s(n17536), .op(n16422) );
  mux2_1 U18398 ( .ip1(\x[64][10] ), .ip2(n17356), .s(n17536), .op(n16421) );
  buf_1 U18399 ( .ip(n17536), .op(n17535) );
  mux2_1 U18400 ( .ip1(\x[64][9] ), .ip2(n17357), .s(n17535), .op(n16420) );
  mux2_1 U18401 ( .ip1(\x[64][8] ), .ip2(n17358), .s(n17536), .op(n16419) );
  mux2_1 U18402 ( .ip1(\x[64][7] ), .ip2(n17359), .s(n17535), .op(n16418) );
  mux2_1 U18403 ( .ip1(\x[64][6] ), .ip2(n17360), .s(n17536), .op(n16417) );
  mux2_1 U18404 ( .ip1(\x[64][5] ), .ip2(n17361), .s(n17535), .op(n16416) );
  mux2_1 U18405 ( .ip1(\x[64][4] ), .ip2(n17362), .s(n17536), .op(n16415) );
  mux2_1 U18406 ( .ip1(\x[64][3] ), .ip2(n17363), .s(n17535), .op(n16414) );
  mux2_1 U18407 ( .ip1(\x[64][2] ), .ip2(n17364), .s(n17535), .op(n16413) );
  mux2_1 U18408 ( .ip1(\x[64][1] ), .ip2(n17365), .s(n17535), .op(n16412) );
  mux2_1 U18409 ( .ip1(\x[64][0] ), .ip2(n17366), .s(n17535), .op(n16411) );
  inv_1 U18410 ( .ip(address[6]), .op(n17371) );
  nand4_1 U18411 ( .ip1(address[4]), .ip2(we), .ip3(address[5]), .ip4(n17371), 
        .op(n17367) );
  nor2_1 U18412 ( .ip1(n17373), .ip2(n17367), .op(n17538) );
  mux2_1 U18413 ( .ip1(\x[63][15] ), .ip2(n17351), .s(n17538), .op(n16410) );
  mux2_1 U18414 ( .ip1(\x[63][14] ), .ip2(n17352), .s(n17538), .op(n16409) );
  mux2_1 U18415 ( .ip1(\x[63][13] ), .ip2(n17353), .s(n17538), .op(n16408) );
  mux2_1 U18416 ( .ip1(\x[63][12] ), .ip2(n17354), .s(n17538), .op(n16407) );
  mux2_1 U18417 ( .ip1(\x[63][11] ), .ip2(n17355), .s(n17538), .op(n16406) );
  mux2_1 U18418 ( .ip1(\x[63][10] ), .ip2(n17356), .s(n17538), .op(n16405) );
  buf_1 U18419 ( .ip(n17538), .op(n17537) );
  mux2_1 U18420 ( .ip1(\x[63][9] ), .ip2(n17357), .s(n17537), .op(n16404) );
  mux2_1 U18421 ( .ip1(\x[63][8] ), .ip2(n17358), .s(n17538), .op(n16403) );
  mux2_1 U18422 ( .ip1(\x[63][7] ), .ip2(n17359), .s(n17537), .op(n16402) );
  mux2_1 U18423 ( .ip1(\x[63][6] ), .ip2(n17360), .s(n17538), .op(n16401) );
  mux2_1 U18424 ( .ip1(\x[63][5] ), .ip2(n17361), .s(n17537), .op(n16400) );
  mux2_1 U18425 ( .ip1(\x[63][4] ), .ip2(n17362), .s(n17538), .op(n16399) );
  mux2_1 U18426 ( .ip1(\x[63][3] ), .ip2(n17363), .s(n17537), .op(n16398) );
  mux2_1 U18427 ( .ip1(\x[63][2] ), .ip2(n17364), .s(n17537), .op(n16397) );
  mux2_1 U18428 ( .ip1(\x[63][1] ), .ip2(n17365), .s(n17537), .op(n16396) );
  mux2_1 U18429 ( .ip1(\x[63][0] ), .ip2(n17366), .s(n17537), .op(n16395) );
  nor2_1 U18430 ( .ip1(n17374), .ip2(n17367), .op(n17540) );
  mux2_1 U18431 ( .ip1(\x[62][15] ), .ip2(n17351), .s(n17540), .op(n16394) );
  mux2_1 U18432 ( .ip1(\x[62][14] ), .ip2(n17352), .s(n17540), .op(n16393) );
  mux2_1 U18433 ( .ip1(\x[62][13] ), .ip2(n17353), .s(n17540), .op(n16392) );
  mux2_1 U18434 ( .ip1(\x[62][12] ), .ip2(n17354), .s(n17540), .op(n16391) );
  mux2_1 U18435 ( .ip1(\x[62][11] ), .ip2(n17355), .s(n17540), .op(n16390) );
  mux2_1 U18436 ( .ip1(\x[62][10] ), .ip2(n17356), .s(n17540), .op(n16389) );
  buf_1 U18437 ( .ip(n17540), .op(n17539) );
  mux2_1 U18438 ( .ip1(\x[62][9] ), .ip2(n17357), .s(n17539), .op(n16388) );
  mux2_1 U18439 ( .ip1(\x[62][8] ), .ip2(n17358), .s(n17540), .op(n16387) );
  mux2_1 U18440 ( .ip1(\x[62][7] ), .ip2(n17359), .s(n17539), .op(n16386) );
  mux2_1 U18441 ( .ip1(\x[62][6] ), .ip2(n17360), .s(n17540), .op(n16385) );
  mux2_1 U18442 ( .ip1(\x[62][5] ), .ip2(n17361), .s(n17539), .op(n16384) );
  mux2_1 U18443 ( .ip1(\x[62][4] ), .ip2(n17362), .s(n17540), .op(n16383) );
  mux2_1 U18444 ( .ip1(\x[62][3] ), .ip2(n17363), .s(n17539), .op(n16382) );
  mux2_1 U18445 ( .ip1(\x[62][2] ), .ip2(n17364), .s(n17539), .op(n16381) );
  mux2_1 U18446 ( .ip1(\x[62][1] ), .ip2(n17365), .s(n17539), .op(n16380) );
  mux2_1 U18447 ( .ip1(\x[62][0] ), .ip2(n17366), .s(n17539), .op(n16379) );
  nor2_1 U18448 ( .ip1(n17375), .ip2(n17367), .op(n17557) );
  mux2_1 U18449 ( .ip1(\x[61][15] ), .ip2(n17351), .s(n17557), .op(n16378) );
  mux2_1 U18450 ( .ip1(\x[61][14] ), .ip2(n17352), .s(n17557), .op(n16377) );
  mux2_1 U18451 ( .ip1(\x[61][13] ), .ip2(n17353), .s(n17557), .op(n16376) );
  mux2_1 U18452 ( .ip1(\x[61][12] ), .ip2(n17354), .s(n17557), .op(n16375) );
  mux2_1 U18453 ( .ip1(\x[61][11] ), .ip2(n17355), .s(n17557), .op(n16374) );
  mux2_1 U18454 ( .ip1(\x[61][10] ), .ip2(n17356), .s(n17557), .op(n16373) );
  buf_1 U18455 ( .ip(n17557), .op(n17550) );
  mux2_1 U18456 ( .ip1(\x[61][9] ), .ip2(n17357), .s(n17550), .op(n16372) );
  mux2_1 U18457 ( .ip1(\x[61][8] ), .ip2(n17358), .s(n17557), .op(n16371) );
  mux2_1 U18458 ( .ip1(\x[61][7] ), .ip2(n17359), .s(n17550), .op(n16370) );
  mux2_1 U18459 ( .ip1(\x[61][6] ), .ip2(n17360), .s(n17557), .op(n16369) );
  mux2_1 U18460 ( .ip1(\x[61][5] ), .ip2(n17361), .s(n17550), .op(n16368) );
  mux2_1 U18461 ( .ip1(\x[61][4] ), .ip2(n17362), .s(n17557), .op(n16367) );
  mux2_1 U18462 ( .ip1(\x[61][3] ), .ip2(n17363), .s(n17550), .op(n16366) );
  mux2_1 U18463 ( .ip1(\x[61][2] ), .ip2(n17364), .s(n17550), .op(n16365) );
  mux2_1 U18464 ( .ip1(\x[61][1] ), .ip2(n17365), .s(n17550), .op(n16364) );
  mux2_1 U18465 ( .ip1(\x[61][0] ), .ip2(n17366), .s(n17550), .op(n16363) );
  nor2_1 U18466 ( .ip1(n17392), .ip2(n17367), .op(n17560) );
  mux2_1 U18467 ( .ip1(\x[60][15] ), .ip2(n17351), .s(n17560), .op(n16362) );
  mux2_1 U18468 ( .ip1(\x[60][14] ), .ip2(n17352), .s(n17560), .op(n16361) );
  mux2_1 U18469 ( .ip1(\x[60][13] ), .ip2(n17353), .s(n17560), .op(n16360) );
  mux2_1 U18470 ( .ip1(\x[60][12] ), .ip2(n17354), .s(n17560), .op(n16359) );
  mux2_1 U18471 ( .ip1(\x[60][11] ), .ip2(n17355), .s(n17560), .op(n16358) );
  mux2_1 U18472 ( .ip1(\x[60][10] ), .ip2(n17356), .s(n17560), .op(n16357) );
  buf_1 U18473 ( .ip(n17560), .op(n17559) );
  mux2_1 U18474 ( .ip1(\x[60][9] ), .ip2(n17357), .s(n17559), .op(n16356) );
  mux2_1 U18475 ( .ip1(\x[60][8] ), .ip2(n17358), .s(n17560), .op(n16355) );
  mux2_1 U18476 ( .ip1(\x[60][7] ), .ip2(n17359), .s(n17559), .op(n16354) );
  mux2_1 U18477 ( .ip1(\x[60][6] ), .ip2(n17360), .s(n17560), .op(n16353) );
  mux2_1 U18478 ( .ip1(\x[60][5] ), .ip2(n17361), .s(n17559), .op(n16352) );
  mux2_1 U18479 ( .ip1(\x[60][4] ), .ip2(n17362), .s(n17560), .op(n16351) );
  mux2_1 U18480 ( .ip1(\x[60][3] ), .ip2(n17363), .s(n17559), .op(n16350) );
  mux2_1 U18481 ( .ip1(\x[60][2] ), .ip2(n17364), .s(n17559), .op(n16349) );
  mux2_1 U18482 ( .ip1(\x[60][1] ), .ip2(n17365), .s(n17559), .op(n16348) );
  mux2_1 U18483 ( .ip1(\x[60][0] ), .ip2(n17366), .s(n17559), .op(n16347) );
  nor2_1 U18484 ( .ip1(n17393), .ip2(n17367), .op(n17562) );
  mux2_1 U18485 ( .ip1(\x[59][15] ), .ip2(n17351), .s(n17562), .op(n16346) );
  mux2_1 U18486 ( .ip1(\x[59][14] ), .ip2(n17352), .s(n17562), .op(n16345) );
  mux2_1 U18487 ( .ip1(\x[59][13] ), .ip2(n17353), .s(n17562), .op(n16344) );
  mux2_1 U18488 ( .ip1(\x[59][12] ), .ip2(n17354), .s(n17562), .op(n16343) );
  mux2_1 U18489 ( .ip1(\x[59][11] ), .ip2(n17355), .s(n17562), .op(n16342) );
  mux2_1 U18490 ( .ip1(\x[59][10] ), .ip2(n17356), .s(n17562), .op(n16341) );
  buf_1 U18491 ( .ip(n17562), .op(n17561) );
  mux2_1 U18492 ( .ip1(\x[59][9] ), .ip2(n17357), .s(n17561), .op(n16340) );
  mux2_1 U18493 ( .ip1(\x[59][8] ), .ip2(n17358), .s(n17562), .op(n16339) );
  mux2_1 U18494 ( .ip1(\x[59][7] ), .ip2(n17359), .s(n17561), .op(n16338) );
  mux2_1 U18495 ( .ip1(\x[59][6] ), .ip2(n17360), .s(n17562), .op(n16337) );
  mux2_1 U18496 ( .ip1(\x[59][5] ), .ip2(n17361), .s(n17561), .op(n16336) );
  mux2_1 U18497 ( .ip1(\x[59][4] ), .ip2(n17362), .s(n17562), .op(n16335) );
  mux2_1 U18498 ( .ip1(\x[59][3] ), .ip2(n17363), .s(n17561), .op(n16334) );
  mux2_1 U18499 ( .ip1(\x[59][2] ), .ip2(n17364), .s(n17561), .op(n16333) );
  mux2_1 U18500 ( .ip1(\x[59][1] ), .ip2(n17365), .s(n17561), .op(n16332) );
  mux2_1 U18501 ( .ip1(\x[59][0] ), .ip2(n17366), .s(n17561), .op(n16331) );
  nor2_1 U18502 ( .ip1(n17394), .ip2(n17367), .op(n17564) );
  mux2_1 U18503 ( .ip1(\x[58][15] ), .ip2(n17351), .s(n17564), .op(n16330) );
  mux2_1 U18504 ( .ip1(\x[58][14] ), .ip2(n17352), .s(n17564), .op(n16329) );
  mux2_1 U18505 ( .ip1(\x[58][13] ), .ip2(n17353), .s(n17564), .op(n16328) );
  mux2_1 U18506 ( .ip1(\x[58][12] ), .ip2(n17354), .s(n17564), .op(n16327) );
  mux2_1 U18507 ( .ip1(\x[58][11] ), .ip2(n17355), .s(n17564), .op(n16326) );
  mux2_1 U18508 ( .ip1(\x[58][10] ), .ip2(n17356), .s(n17564), .op(n16325) );
  buf_1 U18509 ( .ip(n17564), .op(n17563) );
  mux2_1 U18510 ( .ip1(\x[58][9] ), .ip2(n17357), .s(n17563), .op(n16324) );
  mux2_1 U18511 ( .ip1(\x[58][8] ), .ip2(n17358), .s(n17564), .op(n16323) );
  mux2_1 U18512 ( .ip1(\x[58][7] ), .ip2(n17359), .s(n17563), .op(n16322) );
  mux2_1 U18513 ( .ip1(\x[58][6] ), .ip2(n17360), .s(n17564), .op(n16321) );
  mux2_1 U18514 ( .ip1(\x[58][5] ), .ip2(n17361), .s(n17563), .op(n16320) );
  mux2_1 U18515 ( .ip1(\x[58][4] ), .ip2(n17362), .s(n17564), .op(n16319) );
  mux2_1 U18516 ( .ip1(\x[58][3] ), .ip2(n17363), .s(n17563), .op(n16318) );
  mux2_1 U18517 ( .ip1(\x[58][2] ), .ip2(n17364), .s(n17563), .op(n16317) );
  mux2_1 U18518 ( .ip1(\x[58][1] ), .ip2(n17365), .s(n17563), .op(n16316) );
  mux2_1 U18519 ( .ip1(\x[58][0] ), .ip2(n17366), .s(n17563), .op(n16315) );
  nor2_1 U18520 ( .ip1(n17395), .ip2(n17367), .op(n17566) );
  mux2_1 U18521 ( .ip1(\x[57][15] ), .ip2(n17351), .s(n17566), .op(n16314) );
  mux2_1 U18522 ( .ip1(\x[57][14] ), .ip2(n17352), .s(n17566), .op(n16313) );
  mux2_1 U18523 ( .ip1(\x[57][13] ), .ip2(n17353), .s(n17566), .op(n16312) );
  mux2_1 U18524 ( .ip1(\x[57][12] ), .ip2(n17354), .s(n17566), .op(n16311) );
  mux2_1 U18525 ( .ip1(\x[57][11] ), .ip2(n17355), .s(n17566), .op(n16310) );
  mux2_1 U18526 ( .ip1(\x[57][10] ), .ip2(n17356), .s(n17566), .op(n16309) );
  buf_1 U18527 ( .ip(n17566), .op(n17565) );
  mux2_1 U18528 ( .ip1(\x[57][9] ), .ip2(n17357), .s(n17565), .op(n16308) );
  mux2_1 U18529 ( .ip1(\x[57][8] ), .ip2(n17358), .s(n17566), .op(n16307) );
  mux2_1 U18530 ( .ip1(\x[57][7] ), .ip2(n17359), .s(n17565), .op(n16306) );
  mux2_1 U18531 ( .ip1(\x[57][6] ), .ip2(n17360), .s(n17566), .op(n16305) );
  mux2_1 U18532 ( .ip1(\x[57][5] ), .ip2(n17361), .s(n17565), .op(n16304) );
  mux2_1 U18533 ( .ip1(\x[57][4] ), .ip2(n17362), .s(n17566), .op(n16303) );
  mux2_1 U18534 ( .ip1(\x[57][3] ), .ip2(n17363), .s(n17565), .op(n16302) );
  mux2_1 U18535 ( .ip1(\x[57][2] ), .ip2(n17364), .s(n17565), .op(n16301) );
  mux2_1 U18536 ( .ip1(\x[57][1] ), .ip2(n17365), .s(n17565), .op(n16300) );
  mux2_1 U18537 ( .ip1(\x[57][0] ), .ip2(n17366), .s(n17565), .op(n16299) );
  nor2_1 U18538 ( .ip1(n17396), .ip2(n17367), .op(n17568) );
  mux2_1 U18539 ( .ip1(\x[56][15] ), .ip2(n17351), .s(n17568), .op(n16298) );
  mux2_1 U18540 ( .ip1(\x[56][14] ), .ip2(n17352), .s(n17568), .op(n16297) );
  mux2_1 U18541 ( .ip1(\x[56][13] ), .ip2(n17353), .s(n17568), .op(n16296) );
  mux2_1 U18542 ( .ip1(\x[56][12] ), .ip2(n17354), .s(n17568), .op(n16295) );
  mux2_1 U18543 ( .ip1(\x[56][11] ), .ip2(n17355), .s(n17568), .op(n16294) );
  mux2_1 U18544 ( .ip1(\x[56][10] ), .ip2(n17356), .s(n17568), .op(n16293) );
  buf_1 U18545 ( .ip(n17568), .op(n17567) );
  mux2_1 U18546 ( .ip1(\x[56][9] ), .ip2(n17357), .s(n17567), .op(n16292) );
  mux2_1 U18547 ( .ip1(\x[56][8] ), .ip2(n17358), .s(n17568), .op(n16291) );
  mux2_1 U18548 ( .ip1(\x[56][7] ), .ip2(n17359), .s(n17567), .op(n16290) );
  mux2_1 U18549 ( .ip1(\x[56][6] ), .ip2(n17360), .s(n17568), .op(n16289) );
  mux2_1 U18550 ( .ip1(\x[56][5] ), .ip2(n17361), .s(n17567), .op(n16288) );
  mux2_1 U18551 ( .ip1(\x[56][4] ), .ip2(n17362), .s(n17568), .op(n16287) );
  mux2_1 U18552 ( .ip1(\x[56][3] ), .ip2(n17363), .s(n17567), .op(n16286) );
  mux2_1 U18553 ( .ip1(\x[56][2] ), .ip2(n17364), .s(n17567), .op(n16285) );
  mux2_1 U18554 ( .ip1(\x[56][1] ), .ip2(n17365), .s(n17567), .op(n16284) );
  mux2_1 U18555 ( .ip1(\x[56][0] ), .ip2(n17366), .s(n17567), .op(n16283) );
  nor2_1 U18556 ( .ip1(n17397), .ip2(n17367), .op(n17570) );
  mux2_1 U18557 ( .ip1(\x[55][15] ), .ip2(n17351), .s(n17570), .op(n16282) );
  mux2_1 U18558 ( .ip1(\x[55][14] ), .ip2(n17352), .s(n17570), .op(n16281) );
  mux2_1 U18559 ( .ip1(\x[55][13] ), .ip2(n17353), .s(n17570), .op(n16280) );
  mux2_1 U18560 ( .ip1(\x[55][12] ), .ip2(n17354), .s(n17570), .op(n16279) );
  mux2_1 U18561 ( .ip1(\x[55][11] ), .ip2(n17355), .s(n17570), .op(n16278) );
  mux2_1 U18562 ( .ip1(\x[55][10] ), .ip2(n17356), .s(n17570), .op(n16277) );
  buf_1 U18563 ( .ip(n17570), .op(n17569) );
  mux2_1 U18564 ( .ip1(\x[55][9] ), .ip2(n17357), .s(n17569), .op(n16276) );
  mux2_1 U18565 ( .ip1(\x[55][8] ), .ip2(n17358), .s(n17570), .op(n16275) );
  mux2_1 U18566 ( .ip1(\x[55][7] ), .ip2(n17359), .s(n17569), .op(n16274) );
  mux2_1 U18567 ( .ip1(\x[55][6] ), .ip2(n17360), .s(n17570), .op(n16273) );
  mux2_1 U18568 ( .ip1(\x[55][5] ), .ip2(n17361), .s(n17569), .op(n16272) );
  mux2_1 U18569 ( .ip1(\x[55][4] ), .ip2(n17362), .s(n17570), .op(n16271) );
  mux2_1 U18570 ( .ip1(\x[55][3] ), .ip2(n17363), .s(n17569), .op(n16270) );
  mux2_1 U18571 ( .ip1(\x[55][2] ), .ip2(n17364), .s(n17569), .op(n16269) );
  mux2_1 U18572 ( .ip1(\x[55][1] ), .ip2(n17365), .s(n17569), .op(n16268) );
  mux2_1 U18573 ( .ip1(\x[55][0] ), .ip2(n17366), .s(n17569), .op(n16267) );
  nor2_1 U18574 ( .ip1(n17398), .ip2(n17367), .op(n17572) );
  mux2_1 U18575 ( .ip1(\x[54][15] ), .ip2(n17351), .s(n17572), .op(n16266) );
  mux2_1 U18576 ( .ip1(\x[54][14] ), .ip2(n17352), .s(n17572), .op(n16265) );
  mux2_1 U18577 ( .ip1(\x[54][13] ), .ip2(n17353), .s(n17572), .op(n16264) );
  mux2_1 U18578 ( .ip1(\x[54][12] ), .ip2(n17354), .s(n17572), .op(n16263) );
  mux2_1 U18579 ( .ip1(\x[54][11] ), .ip2(n17355), .s(n17572), .op(n16262) );
  mux2_1 U18580 ( .ip1(\x[54][10] ), .ip2(n17356), .s(n17572), .op(n16261) );
  buf_1 U18581 ( .ip(n17572), .op(n17571) );
  mux2_1 U18582 ( .ip1(\x[54][9] ), .ip2(n17357), .s(n17571), .op(n16260) );
  mux2_1 U18583 ( .ip1(\x[54][8] ), .ip2(n17358), .s(n17572), .op(n16259) );
  mux2_1 U18584 ( .ip1(\x[54][7] ), .ip2(n17359), .s(n17571), .op(n16258) );
  mux2_1 U18585 ( .ip1(\x[54][6] ), .ip2(n17360), .s(n17572), .op(n16257) );
  mux2_1 U18586 ( .ip1(\x[54][5] ), .ip2(n17361), .s(n17571), .op(n16256) );
  mux2_1 U18587 ( .ip1(\x[54][4] ), .ip2(n17362), .s(n17572), .op(n16255) );
  mux2_1 U18588 ( .ip1(\x[54][3] ), .ip2(n17363), .s(n17571), .op(n16254) );
  mux2_1 U18589 ( .ip1(\x[54][2] ), .ip2(n17364), .s(n17571), .op(n16253) );
  mux2_1 U18590 ( .ip1(\x[54][1] ), .ip2(n17365), .s(n17571), .op(n16252) );
  mux2_1 U18591 ( .ip1(\x[54][0] ), .ip2(n17366), .s(n17571), .op(n16251) );
  nor2_1 U18592 ( .ip1(n17399), .ip2(n17367), .op(n17574) );
  mux2_1 U18593 ( .ip1(\x[53][15] ), .ip2(n17351), .s(n17574), .op(n16250) );
  mux2_1 U18594 ( .ip1(\x[53][14] ), .ip2(n17352), .s(n17574), .op(n16249) );
  mux2_1 U18595 ( .ip1(\x[53][13] ), .ip2(n17353), .s(n17574), .op(n16248) );
  mux2_1 U18596 ( .ip1(\x[53][12] ), .ip2(n17354), .s(n17574), .op(n16247) );
  mux2_1 U18597 ( .ip1(\x[53][11] ), .ip2(n17355), .s(n17574), .op(n16246) );
  mux2_1 U18598 ( .ip1(\x[53][10] ), .ip2(n17356), .s(n17574), .op(n16245) );
  buf_1 U18599 ( .ip(n17574), .op(n17573) );
  mux2_1 U18600 ( .ip1(\x[53][9] ), .ip2(n17357), .s(n17573), .op(n16244) );
  mux2_1 U18601 ( .ip1(\x[53][8] ), .ip2(n17358), .s(n17574), .op(n16243) );
  mux2_1 U18602 ( .ip1(\x[53][7] ), .ip2(n17359), .s(n17573), .op(n16242) );
  mux2_1 U18603 ( .ip1(\x[53][6] ), .ip2(n17360), .s(n17574), .op(n16241) );
  mux2_1 U18604 ( .ip1(\x[53][5] ), .ip2(n17361), .s(n17573), .op(n16240) );
  mux2_1 U18605 ( .ip1(\x[53][4] ), .ip2(n17362), .s(n17574), .op(n16239) );
  mux2_1 U18606 ( .ip1(\x[53][3] ), .ip2(n17363), .s(n17573), .op(n16238) );
  mux2_1 U18607 ( .ip1(\x[53][2] ), .ip2(n17364), .s(n17573), .op(n16237) );
  mux2_1 U18608 ( .ip1(\x[53][1] ), .ip2(n17365), .s(n17573), .op(n16236) );
  mux2_1 U18609 ( .ip1(\x[53][0] ), .ip2(n17366), .s(n17573), .op(n16235) );
  nor2_1 U18610 ( .ip1(n17400), .ip2(n17367), .op(n17576) );
  mux2_1 U18611 ( .ip1(\x[52][15] ), .ip2(n17351), .s(n17576), .op(n16234) );
  mux2_1 U18612 ( .ip1(\x[52][14] ), .ip2(n17352), .s(n17576), .op(n16233) );
  mux2_1 U18613 ( .ip1(\x[52][13] ), .ip2(n17353), .s(n17576), .op(n16232) );
  mux2_1 U18614 ( .ip1(\x[52][12] ), .ip2(n17354), .s(n17576), .op(n16231) );
  mux2_1 U18615 ( .ip1(\x[52][11] ), .ip2(n17355), .s(n17576), .op(n16230) );
  mux2_1 U18616 ( .ip1(\x[52][10] ), .ip2(n17356), .s(n17576), .op(n16229) );
  buf_1 U18617 ( .ip(n17576), .op(n17575) );
  mux2_1 U18618 ( .ip1(\x[52][9] ), .ip2(n17357), .s(n17575), .op(n16228) );
  mux2_1 U18619 ( .ip1(\x[52][8] ), .ip2(n17358), .s(n17576), .op(n16227) );
  mux2_1 U18620 ( .ip1(\x[52][7] ), .ip2(n17359), .s(n17575), .op(n16226) );
  mux2_1 U18621 ( .ip1(\x[52][6] ), .ip2(n17360), .s(n17576), .op(n16225) );
  mux2_1 U18622 ( .ip1(\x[52][5] ), .ip2(n17361), .s(n17575), .op(n16224) );
  mux2_1 U18623 ( .ip1(\x[52][4] ), .ip2(n17362), .s(n17576), .op(n16223) );
  mux2_1 U18624 ( .ip1(\x[52][3] ), .ip2(n17363), .s(n17575), .op(n16222) );
  mux2_1 U18625 ( .ip1(\x[52][2] ), .ip2(n17364), .s(n17575), .op(n16221) );
  mux2_1 U18626 ( .ip1(\x[52][1] ), .ip2(n17365), .s(n17575), .op(n16220) );
  mux2_1 U18627 ( .ip1(\x[52][0] ), .ip2(n17366), .s(n17575), .op(n16219) );
  nor2_1 U18628 ( .ip1(n17401), .ip2(n17367), .op(n17578) );
  mux2_1 U18629 ( .ip1(\x[51][15] ), .ip2(n17351), .s(n17578), .op(n16218) );
  mux2_1 U18630 ( .ip1(\x[51][14] ), .ip2(n17352), .s(n17578), .op(n16217) );
  mux2_1 U18631 ( .ip1(\x[51][13] ), .ip2(n17353), .s(n17578), .op(n16216) );
  mux2_1 U18632 ( .ip1(\x[51][12] ), .ip2(n17354), .s(n17578), .op(n16215) );
  mux2_1 U18633 ( .ip1(\x[51][11] ), .ip2(n17355), .s(n17578), .op(n16214) );
  mux2_1 U18634 ( .ip1(\x[51][10] ), .ip2(n17356), .s(n17578), .op(n16213) );
  buf_1 U18635 ( .ip(n17578), .op(n17577) );
  mux2_1 U18636 ( .ip1(\x[51][9] ), .ip2(n17357), .s(n17577), .op(n16212) );
  mux2_1 U18637 ( .ip1(\x[51][8] ), .ip2(n17358), .s(n17578), .op(n16211) );
  mux2_1 U18638 ( .ip1(\x[51][7] ), .ip2(n17359), .s(n17577), .op(n16210) );
  mux2_1 U18639 ( .ip1(\x[51][6] ), .ip2(n17360), .s(n17578), .op(n16209) );
  mux2_1 U18640 ( .ip1(\x[51][5] ), .ip2(n17361), .s(n17577), .op(n16208) );
  mux2_1 U18641 ( .ip1(\x[51][4] ), .ip2(n17362), .s(n17578), .op(n16207) );
  mux2_1 U18642 ( .ip1(\x[51][3] ), .ip2(n17363), .s(n17577), .op(n16206) );
  mux2_1 U18643 ( .ip1(\x[51][2] ), .ip2(n17364), .s(n17577), .op(n16205) );
  mux2_1 U18644 ( .ip1(\x[51][1] ), .ip2(n17365), .s(n17577), .op(n16204) );
  mux2_1 U18645 ( .ip1(\x[51][0] ), .ip2(n17366), .s(n17577), .op(n16203) );
  nor2_1 U18646 ( .ip1(n17402), .ip2(n17367), .op(n17580) );
  mux2_1 U18647 ( .ip1(\x[50][15] ), .ip2(n17351), .s(n17580), .op(n16202) );
  mux2_1 U18648 ( .ip1(\x[50][14] ), .ip2(n17352), .s(n17580), .op(n16201) );
  mux2_1 U18649 ( .ip1(\x[50][13] ), .ip2(n17353), .s(n17580), .op(n16200) );
  mux2_1 U18650 ( .ip1(\x[50][12] ), .ip2(n17354), .s(n17580), .op(n16199) );
  mux2_1 U18651 ( .ip1(\x[50][11] ), .ip2(n17355), .s(n17580), .op(n16198) );
  mux2_1 U18652 ( .ip1(\x[50][10] ), .ip2(n17356), .s(n17580), .op(n16197) );
  buf_1 U18653 ( .ip(n17580), .op(n17579) );
  mux2_1 U18654 ( .ip1(\x[50][9] ), .ip2(n17357), .s(n17579), .op(n16196) );
  mux2_1 U18655 ( .ip1(\x[50][8] ), .ip2(n17358), .s(n17580), .op(n16195) );
  mux2_1 U18656 ( .ip1(\x[50][7] ), .ip2(n17359), .s(n17579), .op(n16194) );
  mux2_1 U18657 ( .ip1(\x[50][6] ), .ip2(n17360), .s(n17580), .op(n16193) );
  mux2_1 U18658 ( .ip1(\x[50][5] ), .ip2(n17361), .s(n17579), .op(n16192) );
  mux2_1 U18659 ( .ip1(\x[50][4] ), .ip2(n17362), .s(n17580), .op(n16191) );
  mux2_1 U18660 ( .ip1(\x[50][3] ), .ip2(n17363), .s(n17579), .op(n16190) );
  mux2_1 U18661 ( .ip1(\x[50][2] ), .ip2(n17364), .s(n17579), .op(n16189) );
  mux2_1 U18662 ( .ip1(\x[50][1] ), .ip2(n17365), .s(n17579), .op(n16188) );
  mux2_1 U18663 ( .ip1(\x[50][0] ), .ip2(n17366), .s(n17579), .op(n16187) );
  nor2_1 U18664 ( .ip1(n17403), .ip2(n17367), .op(n17582) );
  mux2_1 U18665 ( .ip1(\x[49][15] ), .ip2(d[15]), .s(n17582), .op(n16186) );
  mux2_1 U18666 ( .ip1(\x[49][14] ), .ip2(d[14]), .s(n17582), .op(n16185) );
  mux2_1 U18667 ( .ip1(\x[49][13] ), .ip2(d[13]), .s(n17582), .op(n16184) );
  mux2_1 U18668 ( .ip1(\x[49][12] ), .ip2(d[12]), .s(n17582), .op(n16183) );
  mux2_1 U18669 ( .ip1(\x[49][11] ), .ip2(d[11]), .s(n17582), .op(n16182) );
  mux2_1 U18670 ( .ip1(\x[49][10] ), .ip2(d[10]), .s(n17582), .op(n16181) );
  buf_1 U18671 ( .ip(n17582), .op(n17581) );
  mux2_1 U18672 ( .ip1(\x[49][9] ), .ip2(d[9]), .s(n17581), .op(n16180) );
  mux2_1 U18673 ( .ip1(\x[49][8] ), .ip2(d[8]), .s(n17582), .op(n16179) );
  mux2_1 U18674 ( .ip1(\x[49][7] ), .ip2(d[7]), .s(n17581), .op(n16178) );
  mux2_1 U18675 ( .ip1(\x[49][6] ), .ip2(d[6]), .s(n17582), .op(n16177) );
  mux2_1 U18676 ( .ip1(\x[49][5] ), .ip2(d[5]), .s(n17581), .op(n16176) );
  mux2_1 U18677 ( .ip1(\x[49][4] ), .ip2(d[4]), .s(n17582), .op(n16175) );
  mux2_1 U18678 ( .ip1(\x[49][3] ), .ip2(d[3]), .s(n17581), .op(n16174) );
  mux2_1 U18679 ( .ip1(\x[49][2] ), .ip2(d[2]), .s(n17581), .op(n16173) );
  mux2_1 U18680 ( .ip1(\x[49][1] ), .ip2(d[1]), .s(n17581), .op(n16172) );
  mux2_1 U18681 ( .ip1(\x[49][0] ), .ip2(d[0]), .s(n17581), .op(n16171) );
  buf_1 U18682 ( .ip(d[15]), .op(n17376) );
  nor2_1 U18683 ( .ip1(n17405), .ip2(n17367), .op(n17584) );
  mux2_1 U18684 ( .ip1(\x[48][15] ), .ip2(n17376), .s(n17584), .op(n16170) );
  buf_1 U18685 ( .ip(d[14]), .op(n17377) );
  mux2_1 U18686 ( .ip1(\x[48][14] ), .ip2(n17377), .s(n17584), .op(n16169) );
  buf_1 U18687 ( .ip(d[13]), .op(n17378) );
  mux2_1 U18688 ( .ip1(\x[48][13] ), .ip2(n17378), .s(n17584), .op(n16168) );
  buf_1 U18689 ( .ip(d[12]), .op(n17379) );
  mux2_1 U18690 ( .ip1(\x[48][12] ), .ip2(n17379), .s(n17584), .op(n16167) );
  buf_1 U18691 ( .ip(d[11]), .op(n17380) );
  mux2_1 U18692 ( .ip1(\x[48][11] ), .ip2(n17380), .s(n17584), .op(n16166) );
  buf_1 U18693 ( .ip(d[10]), .op(n17381) );
  mux2_1 U18694 ( .ip1(\x[48][10] ), .ip2(n17381), .s(n17584), .op(n16165) );
  buf_1 U18695 ( .ip(d[9]), .op(n17382) );
  buf_1 U18696 ( .ip(n17584), .op(n17583) );
  mux2_1 U18697 ( .ip1(\x[48][9] ), .ip2(n17382), .s(n17583), .op(n16164) );
  buf_1 U18698 ( .ip(d[8]), .op(n17383) );
  mux2_1 U18699 ( .ip1(\x[48][8] ), .ip2(n17383), .s(n17584), .op(n16163) );
  buf_1 U18700 ( .ip(d[7]), .op(n17384) );
  mux2_1 U18701 ( .ip1(\x[48][7] ), .ip2(n17384), .s(n17583), .op(n16162) );
  buf_1 U18702 ( .ip(d[6]), .op(n17385) );
  mux2_1 U18703 ( .ip1(\x[48][6] ), .ip2(n17385), .s(n17584), .op(n16161) );
  buf_1 U18704 ( .ip(d[5]), .op(n17386) );
  mux2_1 U18705 ( .ip1(\x[48][5] ), .ip2(n17386), .s(n17583), .op(n16160) );
  buf_1 U18706 ( .ip(d[4]), .op(n17387) );
  mux2_1 U18707 ( .ip1(\x[48][4] ), .ip2(n17387), .s(n17584), .op(n16159) );
  buf_1 U18708 ( .ip(d[3]), .op(n17388) );
  mux2_1 U18709 ( .ip1(\x[48][3] ), .ip2(n17388), .s(n17583), .op(n16158) );
  buf_1 U18710 ( .ip(d[2]), .op(n17389) );
  mux2_1 U18711 ( .ip1(\x[48][2] ), .ip2(n17389), .s(n17583), .op(n16157) );
  buf_1 U18712 ( .ip(d[1]), .op(n17390) );
  mux2_1 U18713 ( .ip1(\x[48][1] ), .ip2(n17390), .s(n17583), .op(n16156) );
  buf_1 U18714 ( .ip(d[0]), .op(n17391) );
  mux2_1 U18715 ( .ip1(\x[48][0] ), .ip2(n17391), .s(n17583), .op(n16155) );
  nand3_1 U18716 ( .ip1(address[5]), .ip2(n17372), .ip3(n17371), .op(n17368)
         );
  nor2_1 U18717 ( .ip1(n17373), .ip2(n17368), .op(n17586) );
  mux2_1 U18718 ( .ip1(\x[47][15] ), .ip2(n17376), .s(n17586), .op(n16154) );
  mux2_1 U18719 ( .ip1(\x[47][14] ), .ip2(n17377), .s(n17586), .op(n16153) );
  mux2_1 U18720 ( .ip1(\x[47][13] ), .ip2(n17378), .s(n17586), .op(n16152) );
  mux2_1 U18721 ( .ip1(\x[47][12] ), .ip2(n17379), .s(n17586), .op(n16151) );
  mux2_1 U18722 ( .ip1(\x[47][11] ), .ip2(n17380), .s(n17586), .op(n16150) );
  mux2_1 U18723 ( .ip1(\x[47][10] ), .ip2(n17381), .s(n17586), .op(n16149) );
  buf_1 U18724 ( .ip(n17586), .op(n17585) );
  mux2_1 U18725 ( .ip1(\x[47][9] ), .ip2(n17382), .s(n17585), .op(n16148) );
  mux2_1 U18726 ( .ip1(\x[47][8] ), .ip2(n17383), .s(n17586), .op(n16147) );
  mux2_1 U18727 ( .ip1(\x[47][7] ), .ip2(n17384), .s(n17585), .op(n16146) );
  mux2_1 U18728 ( .ip1(\x[47][6] ), .ip2(n17385), .s(n17586), .op(n16145) );
  mux2_1 U18729 ( .ip1(\x[47][5] ), .ip2(n17386), .s(n17585), .op(n16144) );
  mux2_1 U18730 ( .ip1(\x[47][4] ), .ip2(n17387), .s(n17586), .op(n16143) );
  mux2_1 U18731 ( .ip1(\x[47][3] ), .ip2(n17388), .s(n17585), .op(n16142) );
  mux2_1 U18732 ( .ip1(\x[47][2] ), .ip2(n17389), .s(n17585), .op(n16141) );
  mux2_1 U18733 ( .ip1(\x[47][1] ), .ip2(n17390), .s(n17585), .op(n16140) );
  mux2_1 U18734 ( .ip1(\x[47][0] ), .ip2(n17391), .s(n17585), .op(n16139) );
  nor2_1 U18735 ( .ip1(n17374), .ip2(n17368), .op(n17588) );
  mux2_1 U18736 ( .ip1(\x[46][15] ), .ip2(n17376), .s(n17588), .op(n16138) );
  mux2_1 U18737 ( .ip1(\x[46][14] ), .ip2(n17377), .s(n17588), .op(n16137) );
  mux2_1 U18738 ( .ip1(\x[46][13] ), .ip2(n17378), .s(n17588), .op(n16136) );
  mux2_1 U18739 ( .ip1(\x[46][12] ), .ip2(n17379), .s(n17588), .op(n16135) );
  mux2_1 U18740 ( .ip1(\x[46][11] ), .ip2(n17380), .s(n17588), .op(n16134) );
  mux2_1 U18741 ( .ip1(\x[46][10] ), .ip2(n17381), .s(n17588), .op(n16133) );
  buf_1 U18742 ( .ip(n17588), .op(n17587) );
  mux2_1 U18743 ( .ip1(\x[46][9] ), .ip2(n17382), .s(n17587), .op(n16132) );
  mux2_1 U18744 ( .ip1(\x[46][8] ), .ip2(n17383), .s(n17588), .op(n16131) );
  mux2_1 U18745 ( .ip1(\x[46][7] ), .ip2(n17384), .s(n17587), .op(n16130) );
  mux2_1 U18746 ( .ip1(\x[46][6] ), .ip2(n17385), .s(n17588), .op(n16129) );
  mux2_1 U18747 ( .ip1(\x[46][5] ), .ip2(n17386), .s(n17587), .op(n16128) );
  mux2_1 U18748 ( .ip1(\x[46][4] ), .ip2(n17387), .s(n17588), .op(n16127) );
  mux2_1 U18749 ( .ip1(\x[46][3] ), .ip2(n17388), .s(n17587), .op(n16126) );
  mux2_1 U18750 ( .ip1(\x[46][2] ), .ip2(n17389), .s(n17587), .op(n16125) );
  mux2_1 U18751 ( .ip1(\x[46][1] ), .ip2(n17390), .s(n17587), .op(n16124) );
  mux2_1 U18752 ( .ip1(\x[46][0] ), .ip2(n17391), .s(n17587), .op(n16123) );
  nor2_1 U18753 ( .ip1(n17375), .ip2(n17368), .op(n17590) );
  mux2_1 U18754 ( .ip1(\x[45][15] ), .ip2(n17376), .s(n17590), .op(n16122) );
  mux2_1 U18755 ( .ip1(\x[45][14] ), .ip2(n17377), .s(n17590), .op(n16121) );
  mux2_1 U18756 ( .ip1(\x[45][13] ), .ip2(n17378), .s(n17590), .op(n16120) );
  mux2_1 U18757 ( .ip1(\x[45][12] ), .ip2(n17379), .s(n17590), .op(n16119) );
  mux2_1 U18758 ( .ip1(\x[45][11] ), .ip2(n17380), .s(n17590), .op(n16118) );
  mux2_1 U18759 ( .ip1(\x[45][10] ), .ip2(n17381), .s(n17590), .op(n16117) );
  buf_1 U18760 ( .ip(n17590), .op(n17589) );
  mux2_1 U18761 ( .ip1(\x[45][9] ), .ip2(n17382), .s(n17589), .op(n16116) );
  mux2_1 U18762 ( .ip1(\x[45][8] ), .ip2(n17383), .s(n17590), .op(n16115) );
  mux2_1 U18763 ( .ip1(\x[45][7] ), .ip2(n17384), .s(n17589), .op(n16114) );
  mux2_1 U18764 ( .ip1(\x[45][6] ), .ip2(n17385), .s(n17590), .op(n16113) );
  mux2_1 U18765 ( .ip1(\x[45][5] ), .ip2(n17386), .s(n17589), .op(n16112) );
  mux2_1 U18766 ( .ip1(\x[45][4] ), .ip2(n17387), .s(n17590), .op(n16111) );
  mux2_1 U18767 ( .ip1(\x[45][3] ), .ip2(n17388), .s(n17589), .op(n16110) );
  mux2_1 U18768 ( .ip1(\x[45][2] ), .ip2(n17389), .s(n17589), .op(n16109) );
  mux2_1 U18769 ( .ip1(\x[45][1] ), .ip2(n17390), .s(n17589), .op(n16108) );
  mux2_1 U18770 ( .ip1(\x[45][0] ), .ip2(n17391), .s(n17589), .op(n16107) );
  nor2_1 U18771 ( .ip1(n17392), .ip2(n17368), .op(n17592) );
  mux2_1 U18772 ( .ip1(\x[44][15] ), .ip2(n17376), .s(n17592), .op(n16106) );
  mux2_1 U18773 ( .ip1(\x[44][14] ), .ip2(n17377), .s(n17592), .op(n16105) );
  mux2_1 U18774 ( .ip1(\x[44][13] ), .ip2(n17378), .s(n17592), .op(n16104) );
  mux2_1 U18775 ( .ip1(\x[44][12] ), .ip2(n17379), .s(n17592), .op(n16103) );
  mux2_1 U18776 ( .ip1(\x[44][11] ), .ip2(n17380), .s(n17592), .op(n16102) );
  mux2_1 U18777 ( .ip1(\x[44][10] ), .ip2(n17381), .s(n17592), .op(n16101) );
  buf_1 U18778 ( .ip(n17592), .op(n17591) );
  mux2_1 U18779 ( .ip1(\x[44][9] ), .ip2(n17382), .s(n17591), .op(n16100) );
  mux2_1 U18780 ( .ip1(\x[44][8] ), .ip2(n17383), .s(n17592), .op(n16099) );
  mux2_1 U18781 ( .ip1(\x[44][7] ), .ip2(n17384), .s(n17591), .op(n16098) );
  mux2_1 U18782 ( .ip1(\x[44][6] ), .ip2(n17385), .s(n17592), .op(n16097) );
  mux2_1 U18783 ( .ip1(\x[44][5] ), .ip2(n17386), .s(n17591), .op(n16096) );
  mux2_1 U18784 ( .ip1(\x[44][4] ), .ip2(n17387), .s(n17592), .op(n16095) );
  mux2_1 U18785 ( .ip1(\x[44][3] ), .ip2(n17388), .s(n17591), .op(n16094) );
  mux2_1 U18786 ( .ip1(\x[44][2] ), .ip2(n17389), .s(n17591), .op(n16093) );
  mux2_1 U18787 ( .ip1(\x[44][1] ), .ip2(n17390), .s(n17591), .op(n16092) );
  mux2_1 U18788 ( .ip1(\x[44][0] ), .ip2(n17391), .s(n17591), .op(n16091) );
  nor2_1 U18789 ( .ip1(n17393), .ip2(n17368), .op(n17594) );
  mux2_1 U18790 ( .ip1(\x[43][15] ), .ip2(n17376), .s(n17594), .op(n16090) );
  mux2_1 U18791 ( .ip1(\x[43][14] ), .ip2(n17377), .s(n17594), .op(n16089) );
  mux2_1 U18792 ( .ip1(\x[43][13] ), .ip2(n17378), .s(n17594), .op(n16088) );
  mux2_1 U18793 ( .ip1(\x[43][12] ), .ip2(n17379), .s(n17594), .op(n16087) );
  mux2_1 U18794 ( .ip1(\x[43][11] ), .ip2(n17380), .s(n17594), .op(n16086) );
  mux2_1 U18795 ( .ip1(\x[43][10] ), .ip2(n17381), .s(n17594), .op(n16085) );
  buf_1 U18796 ( .ip(n17594), .op(n17593) );
  mux2_1 U18797 ( .ip1(\x[43][9] ), .ip2(n17382), .s(n17593), .op(n16084) );
  mux2_1 U18798 ( .ip1(\x[43][8] ), .ip2(n17383), .s(n17594), .op(n16083) );
  mux2_1 U18799 ( .ip1(\x[43][7] ), .ip2(n17384), .s(n17593), .op(n16082) );
  mux2_1 U18800 ( .ip1(\x[43][6] ), .ip2(n17385), .s(n17594), .op(n16081) );
  mux2_1 U18801 ( .ip1(\x[43][5] ), .ip2(n17386), .s(n17593), .op(n16080) );
  mux2_1 U18802 ( .ip1(\x[43][4] ), .ip2(n17387), .s(n17594), .op(n16079) );
  mux2_1 U18803 ( .ip1(\x[43][3] ), .ip2(n17388), .s(n17593), .op(n16078) );
  mux2_1 U18804 ( .ip1(\x[43][2] ), .ip2(n17389), .s(n17593), .op(n16077) );
  mux2_1 U18805 ( .ip1(\x[43][1] ), .ip2(n17390), .s(n17593), .op(n16076) );
  mux2_1 U18806 ( .ip1(\x[43][0] ), .ip2(n17391), .s(n17593), .op(n16075) );
  nor2_1 U18807 ( .ip1(n17394), .ip2(n17368), .op(n17596) );
  mux2_1 U18808 ( .ip1(\x[42][15] ), .ip2(n17376), .s(n17596), .op(n16074) );
  mux2_1 U18809 ( .ip1(\x[42][14] ), .ip2(n17377), .s(n17596), .op(n16073) );
  mux2_1 U18810 ( .ip1(\x[42][13] ), .ip2(n17378), .s(n17596), .op(n16072) );
  mux2_1 U18811 ( .ip1(\x[42][12] ), .ip2(n17379), .s(n17596), .op(n16071) );
  mux2_1 U18812 ( .ip1(\x[42][11] ), .ip2(n17380), .s(n17596), .op(n16070) );
  mux2_1 U18813 ( .ip1(\x[42][10] ), .ip2(n17381), .s(n17596), .op(n16069) );
  buf_1 U18814 ( .ip(n17596), .op(n17595) );
  mux2_1 U18815 ( .ip1(\x[42][9] ), .ip2(n17382), .s(n17595), .op(n16068) );
  mux2_1 U18816 ( .ip1(\x[42][8] ), .ip2(n17383), .s(n17596), .op(n16067) );
  mux2_1 U18817 ( .ip1(\x[42][7] ), .ip2(n17384), .s(n17595), .op(n16066) );
  mux2_1 U18818 ( .ip1(\x[42][6] ), .ip2(n17385), .s(n17596), .op(n16065) );
  mux2_1 U18819 ( .ip1(\x[42][5] ), .ip2(n17386), .s(n17595), .op(n16064) );
  mux2_1 U18820 ( .ip1(\x[42][4] ), .ip2(n17387), .s(n17596), .op(n16063) );
  mux2_1 U18821 ( .ip1(\x[42][3] ), .ip2(n17388), .s(n17595), .op(n16062) );
  mux2_1 U18822 ( .ip1(\x[42][2] ), .ip2(n17389), .s(n17595), .op(n16061) );
  mux2_1 U18823 ( .ip1(\x[42][1] ), .ip2(n17390), .s(n17595), .op(n16060) );
  mux2_1 U18824 ( .ip1(\x[42][0] ), .ip2(n17391), .s(n17595), .op(n16059) );
  nor2_1 U18825 ( .ip1(n17395), .ip2(n17368), .op(n17598) );
  mux2_1 U18826 ( .ip1(\x[41][15] ), .ip2(n17376), .s(n17598), .op(n16058) );
  mux2_1 U18827 ( .ip1(\x[41][14] ), .ip2(n17377), .s(n17598), .op(n16057) );
  mux2_1 U18828 ( .ip1(\x[41][13] ), .ip2(n17378), .s(n17598), .op(n16056) );
  mux2_1 U18829 ( .ip1(\x[41][12] ), .ip2(n17379), .s(n17598), .op(n16055) );
  mux2_1 U18830 ( .ip1(\x[41][11] ), .ip2(n17380), .s(n17598), .op(n16054) );
  mux2_1 U18831 ( .ip1(\x[41][10] ), .ip2(n17381), .s(n17598), .op(n16053) );
  buf_1 U18832 ( .ip(n17598), .op(n17597) );
  mux2_1 U18833 ( .ip1(\x[41][9] ), .ip2(n17382), .s(n17597), .op(n16052) );
  mux2_1 U18834 ( .ip1(\x[41][8] ), .ip2(n17383), .s(n17598), .op(n16051) );
  mux2_1 U18835 ( .ip1(\x[41][7] ), .ip2(n17384), .s(n17597), .op(n16050) );
  mux2_1 U18836 ( .ip1(\x[41][6] ), .ip2(n17385), .s(n17598), .op(n16049) );
  mux2_1 U18837 ( .ip1(\x[41][5] ), .ip2(n17386), .s(n17597), .op(n16048) );
  mux2_1 U18838 ( .ip1(\x[41][4] ), .ip2(n17387), .s(n17598), .op(n16047) );
  mux2_1 U18839 ( .ip1(\x[41][3] ), .ip2(n17388), .s(n17597), .op(n16046) );
  mux2_1 U18840 ( .ip1(\x[41][2] ), .ip2(n17389), .s(n17597), .op(n16045) );
  mux2_1 U18841 ( .ip1(\x[41][1] ), .ip2(n17390), .s(n17597), .op(n16044) );
  mux2_1 U18842 ( .ip1(\x[41][0] ), .ip2(n17391), .s(n17597), .op(n16043) );
  nor2_1 U18843 ( .ip1(n17396), .ip2(n17368), .op(n17600) );
  mux2_1 U18844 ( .ip1(\x[40][15] ), .ip2(n17376), .s(n17600), .op(n16042) );
  mux2_1 U18845 ( .ip1(\x[40][14] ), .ip2(n17377), .s(n17600), .op(n16041) );
  mux2_1 U18846 ( .ip1(\x[40][13] ), .ip2(n17378), .s(n17600), .op(n16040) );
  mux2_1 U18847 ( .ip1(\x[40][12] ), .ip2(n17379), .s(n17600), .op(n16039) );
  mux2_1 U18848 ( .ip1(\x[40][11] ), .ip2(n17380), .s(n17600), .op(n16038) );
  mux2_1 U18849 ( .ip1(\x[40][10] ), .ip2(n17381), .s(n17600), .op(n16037) );
  buf_1 U18850 ( .ip(n17600), .op(n17599) );
  mux2_1 U18851 ( .ip1(\x[40][9] ), .ip2(n17382), .s(n17599), .op(n16036) );
  mux2_1 U18852 ( .ip1(\x[40][8] ), .ip2(n17383), .s(n17600), .op(n16035) );
  mux2_1 U18853 ( .ip1(\x[40][7] ), .ip2(n17384), .s(n17599), .op(n16034) );
  mux2_1 U18854 ( .ip1(\x[40][6] ), .ip2(n17385), .s(n17600), .op(n16033) );
  mux2_1 U18855 ( .ip1(\x[40][5] ), .ip2(n17386), .s(n17599), .op(n16032) );
  mux2_1 U18856 ( .ip1(\x[40][4] ), .ip2(n17387), .s(n17600), .op(n16031) );
  mux2_1 U18857 ( .ip1(\x[40][3] ), .ip2(n17388), .s(n17599), .op(n16030) );
  mux2_1 U18858 ( .ip1(\x[40][2] ), .ip2(n17389), .s(n17599), .op(n16029) );
  mux2_1 U18859 ( .ip1(\x[40][1] ), .ip2(n17390), .s(n17599), .op(n16028) );
  mux2_1 U18860 ( .ip1(\x[40][0] ), .ip2(n17391), .s(n17599), .op(n16027) );
  nor2_1 U18861 ( .ip1(n17397), .ip2(n17368), .op(n17602) );
  mux2_1 U18862 ( .ip1(\x[39][15] ), .ip2(n17376), .s(n17602), .op(n16026) );
  mux2_1 U18863 ( .ip1(\x[39][14] ), .ip2(n17377), .s(n17602), .op(n16025) );
  mux2_1 U18864 ( .ip1(\x[39][13] ), .ip2(n17378), .s(n17602), .op(n16024) );
  mux2_1 U18865 ( .ip1(\x[39][12] ), .ip2(n17379), .s(n17602), .op(n16023) );
  mux2_1 U18866 ( .ip1(\x[39][11] ), .ip2(n17380), .s(n17602), .op(n16022) );
  mux2_1 U18867 ( .ip1(\x[39][10] ), .ip2(n17381), .s(n17602), .op(n16021) );
  buf_1 U18868 ( .ip(n17602), .op(n17601) );
  mux2_1 U18869 ( .ip1(\x[39][9] ), .ip2(n17382), .s(n17601), .op(n16020) );
  mux2_1 U18870 ( .ip1(\x[39][8] ), .ip2(n17383), .s(n17602), .op(n16019) );
  mux2_1 U18871 ( .ip1(\x[39][7] ), .ip2(n17384), .s(n17601), .op(n16018) );
  mux2_1 U18872 ( .ip1(\x[39][6] ), .ip2(n17385), .s(n17602), .op(n16017) );
  mux2_1 U18873 ( .ip1(\x[39][5] ), .ip2(n17386), .s(n17601), .op(n16016) );
  mux2_1 U18874 ( .ip1(\x[39][4] ), .ip2(n17387), .s(n17602), .op(n16015) );
  mux2_1 U18875 ( .ip1(\x[39][3] ), .ip2(n17388), .s(n17601), .op(n16014) );
  mux2_1 U18876 ( .ip1(\x[39][2] ), .ip2(n17389), .s(n17601), .op(n16013) );
  mux2_1 U18877 ( .ip1(\x[39][1] ), .ip2(n17390), .s(n17601), .op(n16012) );
  mux2_1 U18878 ( .ip1(\x[39][0] ), .ip2(n17391), .s(n17601), .op(n16011) );
  nor2_1 U18879 ( .ip1(n17398), .ip2(n17368), .op(n17604) );
  mux2_1 U18880 ( .ip1(\x[38][15] ), .ip2(n17376), .s(n17604), .op(n16010) );
  mux2_1 U18881 ( .ip1(\x[38][14] ), .ip2(n17377), .s(n17604), .op(n16009) );
  mux2_1 U18882 ( .ip1(\x[38][13] ), .ip2(n17378), .s(n17604), .op(n16008) );
  mux2_1 U18883 ( .ip1(\x[38][12] ), .ip2(n17379), .s(n17604), .op(n16007) );
  mux2_1 U18884 ( .ip1(\x[38][11] ), .ip2(n17380), .s(n17604), .op(n16006) );
  mux2_1 U18885 ( .ip1(\x[38][10] ), .ip2(n17381), .s(n17604), .op(n16005) );
  buf_1 U18886 ( .ip(n17604), .op(n17603) );
  mux2_1 U18887 ( .ip1(\x[38][9] ), .ip2(n17382), .s(n17603), .op(n16004) );
  mux2_1 U18888 ( .ip1(\x[38][8] ), .ip2(n17383), .s(n17604), .op(n16003) );
  mux2_1 U18889 ( .ip1(\x[38][7] ), .ip2(n17384), .s(n17603), .op(n16002) );
  mux2_1 U18890 ( .ip1(\x[38][6] ), .ip2(n17385), .s(n17604), .op(n16001) );
  mux2_1 U18891 ( .ip1(\x[38][5] ), .ip2(n17386), .s(n17603), .op(n16000) );
  mux2_1 U18892 ( .ip1(\x[38][4] ), .ip2(n17387), .s(n17604), .op(n15999) );
  mux2_1 U18893 ( .ip1(\x[38][3] ), .ip2(n17388), .s(n17603), .op(n15998) );
  mux2_1 U18894 ( .ip1(\x[38][2] ), .ip2(n17389), .s(n17603), .op(n15997) );
  mux2_1 U18895 ( .ip1(\x[38][1] ), .ip2(n17390), .s(n17603), .op(n15996) );
  mux2_1 U18896 ( .ip1(\x[38][0] ), .ip2(n17391), .s(n17603), .op(n15995) );
  nor2_1 U18897 ( .ip1(n17399), .ip2(n17368), .op(n17606) );
  mux2_1 U18898 ( .ip1(\x[37][15] ), .ip2(n17376), .s(n17606), .op(n15994) );
  mux2_1 U18899 ( .ip1(\x[37][14] ), .ip2(n17377), .s(n17606), .op(n15993) );
  mux2_1 U18900 ( .ip1(\x[37][13] ), .ip2(n17378), .s(n17606), .op(n15992) );
  mux2_1 U18901 ( .ip1(\x[37][12] ), .ip2(n17379), .s(n17606), .op(n15991) );
  mux2_1 U18902 ( .ip1(\x[37][11] ), .ip2(n17380), .s(n17606), .op(n15990) );
  mux2_1 U18903 ( .ip1(\x[37][10] ), .ip2(n17381), .s(n17606), .op(n15989) );
  buf_1 U18904 ( .ip(n17606), .op(n17605) );
  mux2_1 U18905 ( .ip1(\x[37][9] ), .ip2(n17382), .s(n17605), .op(n15988) );
  mux2_1 U18906 ( .ip1(\x[37][8] ), .ip2(n17383), .s(n17606), .op(n15987) );
  mux2_1 U18907 ( .ip1(\x[37][7] ), .ip2(n17384), .s(n17605), .op(n15986) );
  mux2_1 U18908 ( .ip1(\x[37][6] ), .ip2(n17385), .s(n17606), .op(n15985) );
  mux2_1 U18909 ( .ip1(\x[37][5] ), .ip2(n17386), .s(n17605), .op(n15984) );
  mux2_1 U18910 ( .ip1(\x[37][4] ), .ip2(n17387), .s(n17606), .op(n15983) );
  mux2_1 U18911 ( .ip1(\x[37][3] ), .ip2(n17388), .s(n17605), .op(n15982) );
  mux2_1 U18912 ( .ip1(\x[37][2] ), .ip2(n17389), .s(n17605), .op(n15981) );
  mux2_1 U18913 ( .ip1(\x[37][1] ), .ip2(n17390), .s(n17605), .op(n15980) );
  mux2_1 U18914 ( .ip1(\x[37][0] ), .ip2(n17391), .s(n17605), .op(n15979) );
  nor2_1 U18915 ( .ip1(n17400), .ip2(n17368), .op(n17608) );
  mux2_1 U18916 ( .ip1(\x[36][15] ), .ip2(n17376), .s(n17608), .op(n15978) );
  mux2_1 U18917 ( .ip1(\x[36][14] ), .ip2(n17377), .s(n17608), .op(n15977) );
  mux2_1 U18918 ( .ip1(\x[36][13] ), .ip2(n17378), .s(n17608), .op(n15976) );
  mux2_1 U18919 ( .ip1(\x[36][12] ), .ip2(n17379), .s(n17608), .op(n15975) );
  mux2_1 U18920 ( .ip1(\x[36][11] ), .ip2(n17380), .s(n17608), .op(n15974) );
  mux2_1 U18921 ( .ip1(\x[36][10] ), .ip2(n17381), .s(n17608), .op(n15973) );
  buf_1 U18922 ( .ip(n17608), .op(n17607) );
  mux2_1 U18923 ( .ip1(\x[36][9] ), .ip2(n17382), .s(n17607), .op(n15972) );
  mux2_1 U18924 ( .ip1(\x[36][8] ), .ip2(n17383), .s(n17608), .op(n15971) );
  mux2_1 U18925 ( .ip1(\x[36][7] ), .ip2(n17384), .s(n17607), .op(n15970) );
  mux2_1 U18926 ( .ip1(\x[36][6] ), .ip2(n17385), .s(n17608), .op(n15969) );
  mux2_1 U18927 ( .ip1(\x[36][5] ), .ip2(n17386), .s(n17607), .op(n15968) );
  mux2_1 U18928 ( .ip1(\x[36][4] ), .ip2(n17387), .s(n17608), .op(n15967) );
  mux2_1 U18929 ( .ip1(\x[36][3] ), .ip2(n17388), .s(n17607), .op(n15966) );
  mux2_1 U18930 ( .ip1(\x[36][2] ), .ip2(n17389), .s(n17607), .op(n15965) );
  mux2_1 U18931 ( .ip1(\x[36][1] ), .ip2(n17390), .s(n17607), .op(n15964) );
  mux2_1 U18932 ( .ip1(\x[36][0] ), .ip2(n17391), .s(n17607), .op(n15963) );
  nor2_1 U18933 ( .ip1(n17401), .ip2(n17368), .op(n17610) );
  mux2_1 U18934 ( .ip1(\x[35][15] ), .ip2(n17376), .s(n17610), .op(n15962) );
  mux2_1 U18935 ( .ip1(\x[35][14] ), .ip2(n17377), .s(n17610), .op(n15961) );
  mux2_1 U18936 ( .ip1(\x[35][13] ), .ip2(n17378), .s(n17610), .op(n15960) );
  mux2_1 U18937 ( .ip1(\x[35][12] ), .ip2(n17379), .s(n17610), .op(n15959) );
  mux2_1 U18938 ( .ip1(\x[35][11] ), .ip2(n17380), .s(n17610), .op(n15958) );
  mux2_1 U18939 ( .ip1(\x[35][10] ), .ip2(n17381), .s(n17610), .op(n15957) );
  buf_1 U18940 ( .ip(n17610), .op(n17609) );
  mux2_1 U18941 ( .ip1(\x[35][9] ), .ip2(n17382), .s(n17609), .op(n15956) );
  mux2_1 U18942 ( .ip1(\x[35][8] ), .ip2(n17383), .s(n17610), .op(n15955) );
  mux2_1 U18943 ( .ip1(\x[35][7] ), .ip2(n17384), .s(n17609), .op(n15954) );
  mux2_1 U18944 ( .ip1(\x[35][6] ), .ip2(n17385), .s(n17610), .op(n15953) );
  mux2_1 U18945 ( .ip1(\x[35][5] ), .ip2(n17386), .s(n17609), .op(n15952) );
  mux2_1 U18946 ( .ip1(\x[35][4] ), .ip2(n17387), .s(n17610), .op(n15951) );
  mux2_1 U18947 ( .ip1(\x[35][3] ), .ip2(n17388), .s(n17609), .op(n15950) );
  mux2_1 U18948 ( .ip1(\x[35][2] ), .ip2(n17389), .s(n17609), .op(n15949) );
  mux2_1 U18949 ( .ip1(\x[35][1] ), .ip2(n17390), .s(n17609), .op(n15948) );
  mux2_1 U18950 ( .ip1(\x[35][0] ), .ip2(n17391), .s(n17609), .op(n15947) );
  nor2_1 U18951 ( .ip1(n17402), .ip2(n17368), .op(n17612) );
  mux2_1 U18952 ( .ip1(\x[34][15] ), .ip2(n17376), .s(n17612), .op(n15946) );
  mux2_1 U18953 ( .ip1(\x[34][14] ), .ip2(n17377), .s(n17612), .op(n15945) );
  mux2_1 U18954 ( .ip1(\x[34][13] ), .ip2(n17378), .s(n17612), .op(n15944) );
  mux2_1 U18955 ( .ip1(\x[34][12] ), .ip2(n17379), .s(n17612), .op(n15943) );
  mux2_1 U18956 ( .ip1(\x[34][11] ), .ip2(n17380), .s(n17612), .op(n15942) );
  mux2_1 U18957 ( .ip1(\x[34][10] ), .ip2(n17381), .s(n17612), .op(n15941) );
  buf_1 U18958 ( .ip(n17612), .op(n17611) );
  mux2_1 U18959 ( .ip1(\x[34][9] ), .ip2(n17382), .s(n17611), .op(n15940) );
  mux2_1 U18960 ( .ip1(\x[34][8] ), .ip2(n17383), .s(n17612), .op(n15939) );
  mux2_1 U18961 ( .ip1(\x[34][7] ), .ip2(n17384), .s(n17611), .op(n15938) );
  mux2_1 U18962 ( .ip1(\x[34][6] ), .ip2(n17385), .s(n17612), .op(n15937) );
  mux2_1 U18963 ( .ip1(\x[34][5] ), .ip2(n17386), .s(n17611), .op(n15936) );
  mux2_1 U18964 ( .ip1(\x[34][4] ), .ip2(n17387), .s(n17612), .op(n15935) );
  mux2_1 U18965 ( .ip1(\x[34][3] ), .ip2(n17388), .s(n17611), .op(n15934) );
  mux2_1 U18966 ( .ip1(\x[34][2] ), .ip2(n17389), .s(n17611), .op(n15933) );
  mux2_1 U18967 ( .ip1(\x[34][1] ), .ip2(n17390), .s(n17611), .op(n15932) );
  mux2_1 U18968 ( .ip1(\x[34][0] ), .ip2(n17391), .s(n17611), .op(n15931) );
  nor2_1 U18969 ( .ip1(n17403), .ip2(n17368), .op(n17614) );
  mux2_1 U18970 ( .ip1(\x[33][15] ), .ip2(n17376), .s(n17614), .op(n15930) );
  mux2_1 U18971 ( .ip1(\x[33][14] ), .ip2(n17377), .s(n17614), .op(n15929) );
  mux2_1 U18972 ( .ip1(\x[33][13] ), .ip2(n17378), .s(n17614), .op(n15928) );
  mux2_1 U18973 ( .ip1(\x[33][12] ), .ip2(n17379), .s(n17614), .op(n15927) );
  mux2_1 U18974 ( .ip1(\x[33][11] ), .ip2(n17380), .s(n17614), .op(n15926) );
  mux2_1 U18975 ( .ip1(\x[33][10] ), .ip2(n17381), .s(n17614), .op(n15925) );
  buf_1 U18976 ( .ip(n17614), .op(n17613) );
  mux2_1 U18977 ( .ip1(\x[33][9] ), .ip2(n17382), .s(n17613), .op(n15924) );
  mux2_1 U18978 ( .ip1(\x[33][8] ), .ip2(n17383), .s(n17614), .op(n15923) );
  mux2_1 U18979 ( .ip1(\x[33][7] ), .ip2(n17384), .s(n17613), .op(n15922) );
  mux2_1 U18980 ( .ip1(\x[33][6] ), .ip2(n17385), .s(n17614), .op(n15921) );
  mux2_1 U18981 ( .ip1(\x[33][5] ), .ip2(n17386), .s(n17613), .op(n15920) );
  mux2_1 U18982 ( .ip1(\x[33][4] ), .ip2(n17387), .s(n17614), .op(n15919) );
  mux2_1 U18983 ( .ip1(\x[33][3] ), .ip2(n17388), .s(n17613), .op(n15918) );
  mux2_1 U18984 ( .ip1(\x[33][2] ), .ip2(n17389), .s(n17613), .op(n15917) );
  mux2_1 U18985 ( .ip1(\x[33][1] ), .ip2(n17390), .s(n17613), .op(n15916) );
  mux2_1 U18986 ( .ip1(\x[33][0] ), .ip2(n17391), .s(n17613), .op(n15915) );
  nor2_1 U18987 ( .ip1(n17405), .ip2(n17368), .op(n17616) );
  mux2_1 U18988 ( .ip1(\x[32][15] ), .ip2(n17376), .s(n17616), .op(n15914) );
  mux2_1 U18989 ( .ip1(\x[32][14] ), .ip2(n17377), .s(n17616), .op(n15913) );
  mux2_1 U18990 ( .ip1(\x[32][13] ), .ip2(n17378), .s(n17616), .op(n15912) );
  mux2_1 U18991 ( .ip1(\x[32][12] ), .ip2(n17379), .s(n17616), .op(n15911) );
  mux2_1 U18992 ( .ip1(\x[32][11] ), .ip2(n17380), .s(n17616), .op(n15910) );
  mux2_1 U18993 ( .ip1(\x[32][10] ), .ip2(n17381), .s(n17616), .op(n15909) );
  buf_1 U18994 ( .ip(n17616), .op(n17615) );
  mux2_1 U18995 ( .ip1(\x[32][9] ), .ip2(n17382), .s(n17615), .op(n15908) );
  mux2_1 U18996 ( .ip1(\x[32][8] ), .ip2(n17383), .s(n17616), .op(n15907) );
  mux2_1 U18997 ( .ip1(\x[32][7] ), .ip2(n17384), .s(n17615), .op(n15906) );
  mux2_1 U18998 ( .ip1(\x[32][6] ), .ip2(n17385), .s(n17616), .op(n15905) );
  mux2_1 U18999 ( .ip1(\x[32][5] ), .ip2(n17386), .s(n17615), .op(n15904) );
  mux2_1 U19000 ( .ip1(\x[32][4] ), .ip2(n17387), .s(n17616), .op(n15903) );
  mux2_1 U19001 ( .ip1(\x[32][3] ), .ip2(n17388), .s(n17615), .op(n15902) );
  mux2_1 U19002 ( .ip1(\x[32][2] ), .ip2(n17389), .s(n17615), .op(n15901) );
  mux2_1 U19003 ( .ip1(\x[32][1] ), .ip2(n17390), .s(n17615), .op(n15900) );
  mux2_1 U19004 ( .ip1(\x[32][0] ), .ip2(n17391), .s(n17615), .op(n15899) );
  nand4_1 U19005 ( .ip1(address[4]), .ip2(we), .ip3(n17371), .ip4(n17370), 
        .op(n17369) );
  nor2_1 U19006 ( .ip1(n17373), .ip2(n17369), .op(n17618) );
  mux2_1 U19007 ( .ip1(\x[31][15] ), .ip2(n17376), .s(n17618), .op(n15898) );
  mux2_1 U19008 ( .ip1(\x[31][14] ), .ip2(n17377), .s(n17618), .op(n15897) );
  mux2_1 U19009 ( .ip1(\x[31][13] ), .ip2(n17378), .s(n17618), .op(n15896) );
  mux2_1 U19010 ( .ip1(\x[31][12] ), .ip2(n17379), .s(n17618), .op(n15895) );
  mux2_1 U19011 ( .ip1(\x[31][11] ), .ip2(n17380), .s(n17618), .op(n15894) );
  mux2_1 U19012 ( .ip1(\x[31][10] ), .ip2(n17381), .s(n17618), .op(n15893) );
  buf_1 U19013 ( .ip(n17618), .op(n17617) );
  mux2_1 U19014 ( .ip1(\x[31][9] ), .ip2(n17382), .s(n17617), .op(n15892) );
  mux2_1 U19015 ( .ip1(\x[31][8] ), .ip2(n17383), .s(n17618), .op(n15891) );
  mux2_1 U19016 ( .ip1(\x[31][7] ), .ip2(n17384), .s(n17617), .op(n15890) );
  mux2_1 U19017 ( .ip1(\x[31][6] ), .ip2(n17385), .s(n17618), .op(n15889) );
  mux2_1 U19018 ( .ip1(\x[31][5] ), .ip2(n17386), .s(n17617), .op(n15888) );
  mux2_1 U19019 ( .ip1(\x[31][4] ), .ip2(n17387), .s(n17618), .op(n15887) );
  mux2_1 U19020 ( .ip1(\x[31][3] ), .ip2(n17388), .s(n17617), .op(n15886) );
  mux2_1 U19021 ( .ip1(\x[31][2] ), .ip2(n17389), .s(n17617), .op(n15885) );
  mux2_1 U19022 ( .ip1(\x[31][1] ), .ip2(n17390), .s(n17617), .op(n15884) );
  mux2_1 U19023 ( .ip1(\x[31][0] ), .ip2(n17391), .s(n17617), .op(n15883) );
  nor2_1 U19024 ( .ip1(n17374), .ip2(n17369), .op(n17620) );
  mux2_1 U19025 ( .ip1(\x[30][15] ), .ip2(n17376), .s(n17620), .op(n15882) );
  mux2_1 U19026 ( .ip1(\x[30][14] ), .ip2(n17377), .s(n17620), .op(n15881) );
  mux2_1 U19027 ( .ip1(\x[30][13] ), .ip2(n17378), .s(n17620), .op(n15880) );
  mux2_1 U19028 ( .ip1(\x[30][12] ), .ip2(n17379), .s(n17620), .op(n15879) );
  mux2_1 U19029 ( .ip1(\x[30][11] ), .ip2(n17380), .s(n17620), .op(n15878) );
  mux2_1 U19030 ( .ip1(\x[30][10] ), .ip2(n17381), .s(n17620), .op(n15877) );
  buf_1 U19031 ( .ip(n17620), .op(n17619) );
  mux2_1 U19032 ( .ip1(\x[30][9] ), .ip2(n17382), .s(n17619), .op(n15876) );
  mux2_1 U19033 ( .ip1(\x[30][8] ), .ip2(n17383), .s(n17620), .op(n15875) );
  mux2_1 U19034 ( .ip1(\x[30][7] ), .ip2(n17384), .s(n17619), .op(n15874) );
  mux2_1 U19035 ( .ip1(\x[30][6] ), .ip2(n17385), .s(n17620), .op(n15873) );
  mux2_1 U19036 ( .ip1(\x[30][5] ), .ip2(n17386), .s(n17619), .op(n15872) );
  mux2_1 U19037 ( .ip1(\x[30][4] ), .ip2(n17387), .s(n17620), .op(n15871) );
  mux2_1 U19038 ( .ip1(\x[30][3] ), .ip2(n17388), .s(n17619), .op(n15870) );
  mux2_1 U19039 ( .ip1(\x[30][2] ), .ip2(n17389), .s(n17619), .op(n15869) );
  mux2_1 U19040 ( .ip1(\x[30][1] ), .ip2(n17390), .s(n17619), .op(n15868) );
  mux2_1 U19041 ( .ip1(\x[30][0] ), .ip2(n17391), .s(n17619), .op(n15867) );
  nor2_1 U19042 ( .ip1(n17375), .ip2(n17369), .op(n17622) );
  mux2_1 U19043 ( .ip1(\x[29][15] ), .ip2(n17376), .s(n17622), .op(n15866) );
  mux2_1 U19044 ( .ip1(\x[29][14] ), .ip2(n17377), .s(n17622), .op(n15865) );
  mux2_1 U19045 ( .ip1(\x[29][13] ), .ip2(n17378), .s(n17622), .op(n15864) );
  mux2_1 U19046 ( .ip1(\x[29][12] ), .ip2(n17379), .s(n17622), .op(n15863) );
  mux2_1 U19047 ( .ip1(\x[29][11] ), .ip2(n17380), .s(n17622), .op(n15862) );
  mux2_1 U19048 ( .ip1(\x[29][10] ), .ip2(n17381), .s(n17622), .op(n15861) );
  buf_1 U19049 ( .ip(n17622), .op(n17621) );
  mux2_1 U19050 ( .ip1(\x[29][9] ), .ip2(n17382), .s(n17621), .op(n15860) );
  mux2_1 U19051 ( .ip1(\x[29][8] ), .ip2(n17383), .s(n17622), .op(n15859) );
  mux2_1 U19052 ( .ip1(\x[29][7] ), .ip2(n17384), .s(n17621), .op(n15858) );
  mux2_1 U19053 ( .ip1(\x[29][6] ), .ip2(n17385), .s(n17622), .op(n15857) );
  mux2_1 U19054 ( .ip1(\x[29][5] ), .ip2(n17386), .s(n17621), .op(n15856) );
  mux2_1 U19055 ( .ip1(\x[29][4] ), .ip2(n17387), .s(n17622), .op(n15855) );
  mux2_1 U19056 ( .ip1(\x[29][3] ), .ip2(n17388), .s(n17621), .op(n15854) );
  mux2_1 U19057 ( .ip1(\x[29][2] ), .ip2(n17389), .s(n17621), .op(n15853) );
  mux2_1 U19058 ( .ip1(\x[29][1] ), .ip2(n17390), .s(n17621), .op(n15852) );
  mux2_1 U19059 ( .ip1(\x[29][0] ), .ip2(n17391), .s(n17621), .op(n15851) );
  nor2_1 U19060 ( .ip1(n17392), .ip2(n17369), .op(n17624) );
  mux2_1 U19061 ( .ip1(\x[28][15] ), .ip2(n17376), .s(n17624), .op(n15850) );
  mux2_1 U19062 ( .ip1(\x[28][14] ), .ip2(n17377), .s(n17624), .op(n15849) );
  mux2_1 U19063 ( .ip1(\x[28][13] ), .ip2(n17378), .s(n17624), .op(n15848) );
  mux2_1 U19064 ( .ip1(\x[28][12] ), .ip2(n17379), .s(n17624), .op(n15847) );
  mux2_1 U19065 ( .ip1(\x[28][11] ), .ip2(n17380), .s(n17624), .op(n15846) );
  mux2_1 U19066 ( .ip1(\x[28][10] ), .ip2(n17381), .s(n17624), .op(n15845) );
  buf_1 U19067 ( .ip(n17624), .op(n17623) );
  mux2_1 U19068 ( .ip1(\x[28][9] ), .ip2(n17382), .s(n17623), .op(n15844) );
  mux2_1 U19069 ( .ip1(\x[28][8] ), .ip2(n17383), .s(n17624), .op(n15843) );
  mux2_1 U19070 ( .ip1(\x[28][7] ), .ip2(n17384), .s(n17623), .op(n15842) );
  mux2_1 U19071 ( .ip1(\x[28][6] ), .ip2(n17385), .s(n17624), .op(n15841) );
  mux2_1 U19072 ( .ip1(\x[28][5] ), .ip2(n17386), .s(n17623), .op(n15840) );
  mux2_1 U19073 ( .ip1(\x[28][4] ), .ip2(n17387), .s(n17624), .op(n15839) );
  mux2_1 U19074 ( .ip1(\x[28][3] ), .ip2(n17388), .s(n17623), .op(n15838) );
  mux2_1 U19075 ( .ip1(\x[28][2] ), .ip2(n17389), .s(n17623), .op(n15837) );
  mux2_1 U19076 ( .ip1(\x[28][1] ), .ip2(n17390), .s(n17623), .op(n15836) );
  mux2_1 U19077 ( .ip1(\x[28][0] ), .ip2(n17391), .s(n17623), .op(n15835) );
  nor2_1 U19078 ( .ip1(n17393), .ip2(n17369), .op(n17626) );
  mux2_1 U19079 ( .ip1(\x[27][15] ), .ip2(n17376), .s(n17626), .op(n15834) );
  mux2_1 U19080 ( .ip1(\x[27][14] ), .ip2(n17377), .s(n17626), .op(n15833) );
  mux2_1 U19081 ( .ip1(\x[27][13] ), .ip2(n17378), .s(n17626), .op(n15832) );
  mux2_1 U19082 ( .ip1(\x[27][12] ), .ip2(n17379), .s(n17626), .op(n15831) );
  mux2_1 U19083 ( .ip1(\x[27][11] ), .ip2(n17380), .s(n17626), .op(n15830) );
  mux2_1 U19084 ( .ip1(\x[27][10] ), .ip2(n17381), .s(n17626), .op(n15829) );
  buf_1 U19085 ( .ip(n17626), .op(n17625) );
  mux2_1 U19086 ( .ip1(\x[27][9] ), .ip2(n17382), .s(n17625), .op(n15828) );
  mux2_1 U19087 ( .ip1(\x[27][8] ), .ip2(n17383), .s(n17626), .op(n15827) );
  mux2_1 U19088 ( .ip1(\x[27][7] ), .ip2(n17384), .s(n17625), .op(n15826) );
  mux2_1 U19089 ( .ip1(\x[27][6] ), .ip2(n17385), .s(n17626), .op(n15825) );
  mux2_1 U19090 ( .ip1(\x[27][5] ), .ip2(n17386), .s(n17625), .op(n15824) );
  mux2_1 U19091 ( .ip1(\x[27][4] ), .ip2(n17387), .s(n17626), .op(n15823) );
  mux2_1 U19092 ( .ip1(\x[27][3] ), .ip2(n17388), .s(n17625), .op(n15822) );
  mux2_1 U19093 ( .ip1(\x[27][2] ), .ip2(n17389), .s(n17625), .op(n15821) );
  mux2_1 U19094 ( .ip1(\x[27][1] ), .ip2(n17390), .s(n17625), .op(n15820) );
  mux2_1 U19095 ( .ip1(\x[27][0] ), .ip2(n17391), .s(n17625), .op(n15819) );
  nor2_1 U19096 ( .ip1(n17394), .ip2(n17369), .op(n17628) );
  mux2_1 U19097 ( .ip1(\x[26][15] ), .ip2(n17376), .s(n17628), .op(n15818) );
  mux2_1 U19098 ( .ip1(\x[26][14] ), .ip2(n17377), .s(n17628), .op(n15817) );
  mux2_1 U19099 ( .ip1(\x[26][13] ), .ip2(n17378), .s(n17628), .op(n15816) );
  mux2_1 U19100 ( .ip1(\x[26][12] ), .ip2(n17379), .s(n17628), .op(n15815) );
  mux2_1 U19101 ( .ip1(\x[26][11] ), .ip2(n17380), .s(n17628), .op(n15814) );
  mux2_1 U19102 ( .ip1(\x[26][10] ), .ip2(n17381), .s(n17628), .op(n15813) );
  buf_1 U19103 ( .ip(n17628), .op(n17627) );
  mux2_1 U19104 ( .ip1(\x[26][9] ), .ip2(n17382), .s(n17627), .op(n15812) );
  mux2_1 U19105 ( .ip1(\x[26][8] ), .ip2(n17383), .s(n17628), .op(n15811) );
  mux2_1 U19106 ( .ip1(\x[26][7] ), .ip2(n17384), .s(n17627), .op(n15810) );
  mux2_1 U19107 ( .ip1(\x[26][6] ), .ip2(n17385), .s(n17628), .op(n15809) );
  mux2_1 U19108 ( .ip1(\x[26][5] ), .ip2(n17386), .s(n17627), .op(n15808) );
  mux2_1 U19109 ( .ip1(\x[26][4] ), .ip2(n17387), .s(n17628), .op(n15807) );
  mux2_1 U19110 ( .ip1(\x[26][3] ), .ip2(n17388), .s(n17627), .op(n15806) );
  mux2_1 U19111 ( .ip1(\x[26][2] ), .ip2(n17389), .s(n17627), .op(n15805) );
  mux2_1 U19112 ( .ip1(\x[26][1] ), .ip2(n17390), .s(n17627), .op(n15804) );
  mux2_1 U19113 ( .ip1(\x[26][0] ), .ip2(n17391), .s(n17627), .op(n15803) );
  nor2_1 U19114 ( .ip1(n17395), .ip2(n17369), .op(n17645) );
  mux2_1 U19115 ( .ip1(\x[25][15] ), .ip2(n17376), .s(n17645), .op(n15802) );
  mux2_1 U19116 ( .ip1(\x[25][14] ), .ip2(n17377), .s(n17645), .op(n15801) );
  mux2_1 U19117 ( .ip1(\x[25][13] ), .ip2(n17378), .s(n17645), .op(n15800) );
  mux2_1 U19118 ( .ip1(\x[25][12] ), .ip2(n17379), .s(n17645), .op(n15799) );
  mux2_1 U19119 ( .ip1(\x[25][11] ), .ip2(n17380), .s(n17645), .op(n15798) );
  mux2_1 U19120 ( .ip1(\x[25][10] ), .ip2(n17381), .s(n17645), .op(n15797) );
  buf_1 U19121 ( .ip(n17645), .op(n17638) );
  mux2_1 U19122 ( .ip1(\x[25][9] ), .ip2(n17382), .s(n17638), .op(n15796) );
  mux2_1 U19123 ( .ip1(\x[25][8] ), .ip2(n17383), .s(n17645), .op(n15795) );
  mux2_1 U19124 ( .ip1(\x[25][7] ), .ip2(n17384), .s(n17638), .op(n15794) );
  mux2_1 U19125 ( .ip1(\x[25][6] ), .ip2(n17385), .s(n17645), .op(n15793) );
  mux2_1 U19126 ( .ip1(\x[25][5] ), .ip2(n17386), .s(n17638), .op(n15792) );
  mux2_1 U19127 ( .ip1(\x[25][4] ), .ip2(n17387), .s(n17645), .op(n15791) );
  mux2_1 U19128 ( .ip1(\x[25][3] ), .ip2(n17388), .s(n17638), .op(n15790) );
  mux2_1 U19129 ( .ip1(\x[25][2] ), .ip2(n17389), .s(n17638), .op(n15789) );
  mux2_1 U19130 ( .ip1(\x[25][1] ), .ip2(n17390), .s(n17638), .op(n15788) );
  mux2_1 U19131 ( .ip1(\x[25][0] ), .ip2(n17391), .s(n17638), .op(n15787) );
  nor2_1 U19132 ( .ip1(n17396), .ip2(n17369), .op(n17648) );
  mux2_1 U19133 ( .ip1(\x[24][15] ), .ip2(n17376), .s(n17648), .op(n15786) );
  mux2_1 U19134 ( .ip1(\x[24][14] ), .ip2(n17377), .s(n17648), .op(n15785) );
  mux2_1 U19135 ( .ip1(\x[24][13] ), .ip2(n17378), .s(n17648), .op(n15784) );
  mux2_1 U19136 ( .ip1(\x[24][12] ), .ip2(n17379), .s(n17648), .op(n15783) );
  mux2_1 U19137 ( .ip1(\x[24][11] ), .ip2(n17380), .s(n17648), .op(n15782) );
  mux2_1 U19138 ( .ip1(\x[24][10] ), .ip2(n17381), .s(n17648), .op(n15781) );
  buf_1 U19139 ( .ip(n17648), .op(n17647) );
  mux2_1 U19140 ( .ip1(\x[24][9] ), .ip2(n17382), .s(n17647), .op(n15780) );
  mux2_1 U19141 ( .ip1(\x[24][8] ), .ip2(n17383), .s(n17648), .op(n15779) );
  mux2_1 U19142 ( .ip1(\x[24][7] ), .ip2(n17384), .s(n17647), .op(n15778) );
  mux2_1 U19143 ( .ip1(\x[24][6] ), .ip2(n17385), .s(n17648), .op(n15777) );
  mux2_1 U19144 ( .ip1(\x[24][5] ), .ip2(n17386), .s(n17647), .op(n15776) );
  mux2_1 U19145 ( .ip1(\x[24][4] ), .ip2(n17387), .s(n17648), .op(n15775) );
  mux2_1 U19146 ( .ip1(\x[24][3] ), .ip2(n17388), .s(n17647), .op(n15774) );
  mux2_1 U19147 ( .ip1(\x[24][2] ), .ip2(n17389), .s(n17647), .op(n15773) );
  mux2_1 U19148 ( .ip1(\x[24][1] ), .ip2(n17390), .s(n17647), .op(n15772) );
  mux2_1 U19149 ( .ip1(\x[24][0] ), .ip2(n17391), .s(n17647), .op(n15771) );
  nor2_1 U19150 ( .ip1(n17397), .ip2(n17369), .op(n17650) );
  mux2_1 U19151 ( .ip1(\x[23][15] ), .ip2(n17376), .s(n17650), .op(n15770) );
  mux2_1 U19152 ( .ip1(\x[23][14] ), .ip2(n17377), .s(n17650), .op(n15769) );
  mux2_1 U19153 ( .ip1(\x[23][13] ), .ip2(n17378), .s(n17650), .op(n15768) );
  mux2_1 U19154 ( .ip1(\x[23][12] ), .ip2(n17379), .s(n17650), .op(n15767) );
  mux2_1 U19155 ( .ip1(\x[23][11] ), .ip2(n17380), .s(n17650), .op(n15766) );
  mux2_1 U19156 ( .ip1(\x[23][10] ), .ip2(n17381), .s(n17650), .op(n15765) );
  buf_1 U19157 ( .ip(n17650), .op(n17649) );
  mux2_1 U19158 ( .ip1(\x[23][9] ), .ip2(n17382), .s(n17649), .op(n15764) );
  mux2_1 U19159 ( .ip1(\x[23][8] ), .ip2(n17383), .s(n17650), .op(n15763) );
  mux2_1 U19160 ( .ip1(\x[23][7] ), .ip2(n17384), .s(n17649), .op(n15762) );
  mux2_1 U19161 ( .ip1(\x[23][6] ), .ip2(n17385), .s(n17650), .op(n15761) );
  mux2_1 U19162 ( .ip1(\x[23][5] ), .ip2(n17386), .s(n17649), .op(n15760) );
  mux2_1 U19163 ( .ip1(\x[23][4] ), .ip2(n17387), .s(n17650), .op(n15759) );
  mux2_1 U19164 ( .ip1(\x[23][3] ), .ip2(n17388), .s(n17649), .op(n15758) );
  mux2_1 U19165 ( .ip1(\x[23][2] ), .ip2(n17389), .s(n17649), .op(n15757) );
  mux2_1 U19166 ( .ip1(\x[23][1] ), .ip2(n17390), .s(n17649), .op(n15756) );
  mux2_1 U19167 ( .ip1(\x[23][0] ), .ip2(n17391), .s(n17649), .op(n15755) );
  nor2_1 U19168 ( .ip1(n17398), .ip2(n17369), .op(n17652) );
  mux2_1 U19169 ( .ip1(\x[22][15] ), .ip2(n17376), .s(n17652), .op(n15754) );
  mux2_1 U19170 ( .ip1(\x[22][14] ), .ip2(n17377), .s(n17652), .op(n15753) );
  mux2_1 U19171 ( .ip1(\x[22][13] ), .ip2(n17378), .s(n17652), .op(n15752) );
  mux2_1 U19172 ( .ip1(\x[22][12] ), .ip2(n17379), .s(n17652), .op(n15751) );
  mux2_1 U19173 ( .ip1(\x[22][11] ), .ip2(n17380), .s(n17652), .op(n15750) );
  mux2_1 U19174 ( .ip1(\x[22][10] ), .ip2(n17381), .s(n17652), .op(n15749) );
  buf_1 U19175 ( .ip(n17652), .op(n17651) );
  mux2_1 U19176 ( .ip1(\x[22][9] ), .ip2(n17382), .s(n17651), .op(n15748) );
  mux2_1 U19177 ( .ip1(\x[22][8] ), .ip2(n17383), .s(n17652), .op(n15747) );
  mux2_1 U19178 ( .ip1(\x[22][7] ), .ip2(n17384), .s(n17651), .op(n15746) );
  mux2_1 U19179 ( .ip1(\x[22][6] ), .ip2(n17385), .s(n17652), .op(n15745) );
  mux2_1 U19180 ( .ip1(\x[22][5] ), .ip2(n17386), .s(n17651), .op(n15744) );
  mux2_1 U19181 ( .ip1(\x[22][4] ), .ip2(n17387), .s(n17652), .op(n15743) );
  mux2_1 U19182 ( .ip1(\x[22][3] ), .ip2(n17388), .s(n17651), .op(n15742) );
  mux2_1 U19183 ( .ip1(\x[22][2] ), .ip2(n17389), .s(n17651), .op(n15741) );
  mux2_1 U19184 ( .ip1(\x[22][1] ), .ip2(n17390), .s(n17651), .op(n15740) );
  mux2_1 U19185 ( .ip1(\x[22][0] ), .ip2(n17391), .s(n17651), .op(n15739) );
  nor2_1 U19186 ( .ip1(n17399), .ip2(n17369), .op(n17654) );
  mux2_1 U19187 ( .ip1(\x[21][15] ), .ip2(n17376), .s(n17654), .op(n15738) );
  mux2_1 U19188 ( .ip1(\x[21][14] ), .ip2(n17377), .s(n17654), .op(n15737) );
  mux2_1 U19189 ( .ip1(\x[21][13] ), .ip2(n17378), .s(n17654), .op(n15736) );
  mux2_1 U19190 ( .ip1(\x[21][12] ), .ip2(n17379), .s(n17654), .op(n15735) );
  mux2_1 U19191 ( .ip1(\x[21][11] ), .ip2(n17380), .s(n17654), .op(n15734) );
  mux2_1 U19192 ( .ip1(\x[21][10] ), .ip2(n17381), .s(n17654), .op(n15733) );
  buf_1 U19193 ( .ip(n17654), .op(n17653) );
  mux2_1 U19194 ( .ip1(\x[21][9] ), .ip2(n17382), .s(n17653), .op(n15732) );
  mux2_1 U19195 ( .ip1(\x[21][8] ), .ip2(n17383), .s(n17654), .op(n15731) );
  mux2_1 U19196 ( .ip1(\x[21][7] ), .ip2(n17384), .s(n17653), .op(n15730) );
  mux2_1 U19197 ( .ip1(\x[21][6] ), .ip2(n17385), .s(n17654), .op(n15729) );
  mux2_1 U19198 ( .ip1(\x[21][5] ), .ip2(n17386), .s(n17653), .op(n15728) );
  mux2_1 U19199 ( .ip1(\x[21][4] ), .ip2(n17387), .s(n17654), .op(n15727) );
  mux2_1 U19200 ( .ip1(\x[21][3] ), .ip2(n17388), .s(n17653), .op(n15726) );
  mux2_1 U19201 ( .ip1(\x[21][2] ), .ip2(n17389), .s(n17653), .op(n15725) );
  mux2_1 U19202 ( .ip1(\x[21][1] ), .ip2(n17390), .s(n17653), .op(n15724) );
  mux2_1 U19203 ( .ip1(\x[21][0] ), .ip2(n17391), .s(n17653), .op(n15723) );
  nor2_1 U19204 ( .ip1(n17400), .ip2(n17369), .op(n17656) );
  mux2_1 U19205 ( .ip1(\x[20][15] ), .ip2(n17376), .s(n17656), .op(n15722) );
  mux2_1 U19206 ( .ip1(\x[20][14] ), .ip2(n17377), .s(n17656), .op(n15721) );
  mux2_1 U19207 ( .ip1(\x[20][13] ), .ip2(n17378), .s(n17656), .op(n15720) );
  mux2_1 U19208 ( .ip1(\x[20][12] ), .ip2(n17379), .s(n17656), .op(n15719) );
  mux2_1 U19209 ( .ip1(\x[20][11] ), .ip2(n17380), .s(n17656), .op(n15718) );
  mux2_1 U19210 ( .ip1(\x[20][10] ), .ip2(n17381), .s(n17656), .op(n15717) );
  buf_1 U19211 ( .ip(n17656), .op(n17655) );
  mux2_1 U19212 ( .ip1(\x[20][9] ), .ip2(n17382), .s(n17655), .op(n15716) );
  mux2_1 U19213 ( .ip1(\x[20][8] ), .ip2(n17383), .s(n17656), .op(n15715) );
  mux2_1 U19214 ( .ip1(\x[20][7] ), .ip2(n17384), .s(n17655), .op(n15714) );
  mux2_1 U19215 ( .ip1(\x[20][6] ), .ip2(n17385), .s(n17656), .op(n15713) );
  mux2_1 U19216 ( .ip1(\x[20][5] ), .ip2(n17386), .s(n17655), .op(n15712) );
  mux2_1 U19217 ( .ip1(\x[20][4] ), .ip2(n17387), .s(n17656), .op(n15711) );
  mux2_1 U19218 ( .ip1(\x[20][3] ), .ip2(n17388), .s(n17655), .op(n15710) );
  mux2_1 U19219 ( .ip1(\x[20][2] ), .ip2(n17389), .s(n17655), .op(n15709) );
  mux2_1 U19220 ( .ip1(\x[20][1] ), .ip2(n17390), .s(n17655), .op(n15708) );
  mux2_1 U19221 ( .ip1(\x[20][0] ), .ip2(n17391), .s(n17655), .op(n15707) );
  nor2_1 U19222 ( .ip1(n17401), .ip2(n17369), .op(n17658) );
  mux2_1 U19223 ( .ip1(\x[19][15] ), .ip2(n17376), .s(n17658), .op(n15706) );
  mux2_1 U19224 ( .ip1(\x[19][14] ), .ip2(n17377), .s(n17658), .op(n15705) );
  mux2_1 U19225 ( .ip1(\x[19][13] ), .ip2(n17378), .s(n17658), .op(n15704) );
  mux2_1 U19226 ( .ip1(\x[19][12] ), .ip2(n17379), .s(n17658), .op(n15703) );
  mux2_1 U19227 ( .ip1(\x[19][11] ), .ip2(n17380), .s(n17658), .op(n15702) );
  mux2_1 U19228 ( .ip1(\x[19][10] ), .ip2(n17381), .s(n17658), .op(n15701) );
  buf_1 U19229 ( .ip(n17658), .op(n17657) );
  mux2_1 U19230 ( .ip1(\x[19][9] ), .ip2(n17382), .s(n17657), .op(n15700) );
  mux2_1 U19231 ( .ip1(\x[19][8] ), .ip2(n17383), .s(n17658), .op(n15699) );
  mux2_1 U19232 ( .ip1(\x[19][7] ), .ip2(n17384), .s(n17657), .op(n15698) );
  mux2_1 U19233 ( .ip1(\x[19][6] ), .ip2(n17385), .s(n17658), .op(n15697) );
  mux2_1 U19234 ( .ip1(\x[19][5] ), .ip2(n17386), .s(n17657), .op(n15696) );
  mux2_1 U19235 ( .ip1(\x[19][4] ), .ip2(n17387), .s(n17658), .op(n15695) );
  mux2_1 U19236 ( .ip1(\x[19][3] ), .ip2(n17388), .s(n17657), .op(n15694) );
  mux2_1 U19237 ( .ip1(\x[19][2] ), .ip2(n17389), .s(n17657), .op(n15693) );
  mux2_1 U19238 ( .ip1(\x[19][1] ), .ip2(n17390), .s(n17657), .op(n15692) );
  mux2_1 U19239 ( .ip1(\x[19][0] ), .ip2(n17391), .s(n17657), .op(n15691) );
  nor2_1 U19240 ( .ip1(n17402), .ip2(n17369), .op(n17660) );
  mux2_1 U19241 ( .ip1(\x[18][15] ), .ip2(n17376), .s(n17660), .op(n15690) );
  mux2_1 U19242 ( .ip1(\x[18][14] ), .ip2(n17377), .s(n17660), .op(n15689) );
  mux2_1 U19243 ( .ip1(\x[18][13] ), .ip2(n17378), .s(n17660), .op(n15688) );
  mux2_1 U19244 ( .ip1(\x[18][12] ), .ip2(n17379), .s(n17660), .op(n15687) );
  mux2_1 U19245 ( .ip1(\x[18][11] ), .ip2(n17380), .s(n17660), .op(n15686) );
  mux2_1 U19246 ( .ip1(\x[18][10] ), .ip2(n17381), .s(n17660), .op(n15685) );
  buf_1 U19247 ( .ip(n17660), .op(n17659) );
  mux2_1 U19248 ( .ip1(\x[18][9] ), .ip2(n17382), .s(n17659), .op(n15684) );
  mux2_1 U19249 ( .ip1(\x[18][8] ), .ip2(n17383), .s(n17660), .op(n15683) );
  mux2_1 U19250 ( .ip1(\x[18][7] ), .ip2(n17384), .s(n17659), .op(n15682) );
  mux2_1 U19251 ( .ip1(\x[18][6] ), .ip2(n17385), .s(n17660), .op(n15681) );
  mux2_1 U19252 ( .ip1(\x[18][5] ), .ip2(n17386), .s(n17659), .op(n15680) );
  mux2_1 U19253 ( .ip1(\x[18][4] ), .ip2(n17387), .s(n17660), .op(n15679) );
  mux2_1 U19254 ( .ip1(\x[18][3] ), .ip2(n17388), .s(n17659), .op(n15678) );
  mux2_1 U19255 ( .ip1(\x[18][2] ), .ip2(n17389), .s(n17659), .op(n15677) );
  mux2_1 U19256 ( .ip1(\x[18][1] ), .ip2(n17390), .s(n17659), .op(n15676) );
  mux2_1 U19257 ( .ip1(\x[18][0] ), .ip2(n17391), .s(n17659), .op(n15675) );
  nor2_1 U19258 ( .ip1(n17403), .ip2(n17369), .op(n17662) );
  mux2_1 U19259 ( .ip1(\x[17][15] ), .ip2(n17376), .s(n17662), .op(n15674) );
  mux2_1 U19260 ( .ip1(\x[17][14] ), .ip2(n17377), .s(n17662), .op(n15673) );
  mux2_1 U19261 ( .ip1(\x[17][13] ), .ip2(n17378), .s(n17662), .op(n15672) );
  mux2_1 U19262 ( .ip1(\x[17][12] ), .ip2(n17379), .s(n17662), .op(n15671) );
  mux2_1 U19263 ( .ip1(\x[17][11] ), .ip2(n17380), .s(n17662), .op(n15670) );
  mux2_1 U19264 ( .ip1(\x[17][10] ), .ip2(n17381), .s(n17662), .op(n15669) );
  buf_1 U19265 ( .ip(n17662), .op(n17661) );
  mux2_1 U19266 ( .ip1(\x[17][9] ), .ip2(n17382), .s(n17661), .op(n15668) );
  mux2_1 U19267 ( .ip1(\x[17][8] ), .ip2(n17383), .s(n17662), .op(n15667) );
  mux2_1 U19268 ( .ip1(\x[17][7] ), .ip2(n17384), .s(n17661), .op(n15666) );
  mux2_1 U19269 ( .ip1(\x[17][6] ), .ip2(n17385), .s(n17662), .op(n15665) );
  mux2_1 U19270 ( .ip1(\x[17][5] ), .ip2(n17386), .s(n17661), .op(n15664) );
  mux2_1 U19271 ( .ip1(\x[17][4] ), .ip2(n17387), .s(n17662), .op(n15663) );
  mux2_1 U19272 ( .ip1(\x[17][3] ), .ip2(n17388), .s(n17661), .op(n15662) );
  mux2_1 U19273 ( .ip1(\x[17][2] ), .ip2(n17389), .s(n17661), .op(n15661) );
  mux2_1 U19274 ( .ip1(\x[17][1] ), .ip2(n17390), .s(n17661), .op(n15660) );
  mux2_1 U19275 ( .ip1(\x[17][0] ), .ip2(n17391), .s(n17661), .op(n15659) );
  nor2_1 U19276 ( .ip1(n17405), .ip2(n17369), .op(n17664) );
  mux2_1 U19277 ( .ip1(\x[16][15] ), .ip2(n17376), .s(n17664), .op(n15658) );
  mux2_1 U19278 ( .ip1(\x[16][14] ), .ip2(n17377), .s(n17664), .op(n15657) );
  mux2_1 U19279 ( .ip1(\x[16][13] ), .ip2(n17378), .s(n17664), .op(n15656) );
  mux2_1 U19280 ( .ip1(\x[16][12] ), .ip2(n17379), .s(n17664), .op(n15655) );
  mux2_1 U19281 ( .ip1(\x[16][11] ), .ip2(n17380), .s(n17664), .op(n15654) );
  mux2_1 U19282 ( .ip1(\x[16][10] ), .ip2(n17381), .s(n17664), .op(n15653) );
  buf_1 U19283 ( .ip(n17664), .op(n17663) );
  mux2_1 U19284 ( .ip1(\x[16][9] ), .ip2(n17382), .s(n17663), .op(n15652) );
  mux2_1 U19285 ( .ip1(\x[16][8] ), .ip2(n17383), .s(n17664), .op(n15651) );
  mux2_1 U19286 ( .ip1(\x[16][7] ), .ip2(n17384), .s(n17663), .op(n15650) );
  mux2_1 U19287 ( .ip1(\x[16][6] ), .ip2(n17385), .s(n17664), .op(n15649) );
  mux2_1 U19288 ( .ip1(\x[16][5] ), .ip2(n17386), .s(n17663), .op(n15648) );
  mux2_1 U19289 ( .ip1(\x[16][4] ), .ip2(n17387), .s(n17664), .op(n15647) );
  mux2_1 U19290 ( .ip1(\x[16][3] ), .ip2(n17388), .s(n17663), .op(n15646) );
  mux2_1 U19291 ( .ip1(\x[16][2] ), .ip2(n17389), .s(n17663), .op(n15645) );
  mux2_1 U19292 ( .ip1(\x[16][1] ), .ip2(n17390), .s(n17663), .op(n15644) );
  mux2_1 U19293 ( .ip1(\x[16][0] ), .ip2(n17391), .s(n17663), .op(n15643) );
  nand3_1 U19294 ( .ip1(n17372), .ip2(n17371), .ip3(n17370), .op(n17404) );
  nor2_1 U19295 ( .ip1(n17373), .ip2(n17404), .op(n17666) );
  mux2_1 U19296 ( .ip1(\x[15][15] ), .ip2(n17376), .s(n17666), .op(n15642) );
  mux2_1 U19297 ( .ip1(\x[15][14] ), .ip2(n17377), .s(n17666), .op(n15641) );
  mux2_1 U19298 ( .ip1(\x[15][13] ), .ip2(n17378), .s(n17666), .op(n15640) );
  mux2_1 U19299 ( .ip1(\x[15][12] ), .ip2(n17379), .s(n17666), .op(n15639) );
  mux2_1 U19300 ( .ip1(\x[15][11] ), .ip2(n17380), .s(n17666), .op(n15638) );
  mux2_1 U19301 ( .ip1(\x[15][10] ), .ip2(n17381), .s(n17666), .op(n15637) );
  buf_1 U19302 ( .ip(n17666), .op(n17665) );
  mux2_1 U19303 ( .ip1(\x[15][9] ), .ip2(n17382), .s(n17665), .op(n15636) );
  mux2_1 U19304 ( .ip1(\x[15][8] ), .ip2(n17383), .s(n17666), .op(n15635) );
  mux2_1 U19305 ( .ip1(\x[15][7] ), .ip2(n17384), .s(n17665), .op(n15634) );
  mux2_1 U19306 ( .ip1(\x[15][6] ), .ip2(n17385), .s(n17666), .op(n15633) );
  mux2_1 U19307 ( .ip1(\x[15][5] ), .ip2(n17386), .s(n17665), .op(n15632) );
  mux2_1 U19308 ( .ip1(\x[15][4] ), .ip2(n17387), .s(n17666), .op(n15631) );
  mux2_1 U19309 ( .ip1(\x[15][3] ), .ip2(n17388), .s(n17665), .op(n15630) );
  mux2_1 U19310 ( .ip1(\x[15][2] ), .ip2(n17389), .s(n17665), .op(n15629) );
  mux2_1 U19311 ( .ip1(\x[15][1] ), .ip2(n17390), .s(n17665), .op(n15628) );
  mux2_1 U19312 ( .ip1(\x[15][0] ), .ip2(n17391), .s(n17665), .op(n15627) );
  nor2_1 U19313 ( .ip1(n17374), .ip2(n17404), .op(n17668) );
  mux2_1 U19314 ( .ip1(\x[14][15] ), .ip2(d[15]), .s(n17668), .op(n15626) );
  mux2_1 U19315 ( .ip1(\x[14][14] ), .ip2(d[14]), .s(n17668), .op(n15625) );
  mux2_1 U19316 ( .ip1(\x[14][13] ), .ip2(d[13]), .s(n17668), .op(n15624) );
  mux2_1 U19317 ( .ip1(\x[14][12] ), .ip2(d[12]), .s(n17668), .op(n15623) );
  mux2_1 U19318 ( .ip1(\x[14][11] ), .ip2(d[11]), .s(n17668), .op(n15622) );
  mux2_1 U19319 ( .ip1(\x[14][10] ), .ip2(d[10]), .s(n17668), .op(n15621) );
  buf_1 U19320 ( .ip(n17668), .op(n17667) );
  mux2_1 U19321 ( .ip1(\x[14][9] ), .ip2(d[9]), .s(n17667), .op(n15620) );
  mux2_1 U19322 ( .ip1(\x[14][8] ), .ip2(d[8]), .s(n17668), .op(n15619) );
  mux2_1 U19323 ( .ip1(\x[14][7] ), .ip2(d[7]), .s(n17667), .op(n15618) );
  mux2_1 U19324 ( .ip1(\x[14][6] ), .ip2(d[6]), .s(n17668), .op(n15617) );
  mux2_1 U19325 ( .ip1(\x[14][5] ), .ip2(d[5]), .s(n17667), .op(n15616) );
  mux2_1 U19326 ( .ip1(\x[14][4] ), .ip2(d[4]), .s(n17668), .op(n15615) );
  mux2_1 U19327 ( .ip1(\x[14][3] ), .ip2(d[3]), .s(n17667), .op(n15614) );
  mux2_1 U19328 ( .ip1(\x[14][2] ), .ip2(d[2]), .s(n17667), .op(n15613) );
  mux2_1 U19329 ( .ip1(\x[14][1] ), .ip2(d[1]), .s(n17667), .op(n15612) );
  mux2_1 U19330 ( .ip1(\x[14][0] ), .ip2(d[0]), .s(n17667), .op(n15611) );
  nor2_1 U19331 ( .ip1(n17375), .ip2(n17404), .op(n17670) );
  mux2_1 U19332 ( .ip1(\x[13][15] ), .ip2(n17376), .s(n17670), .op(n15610) );
  mux2_1 U19333 ( .ip1(\x[13][14] ), .ip2(n17377), .s(n17670), .op(n15609) );
  mux2_1 U19334 ( .ip1(\x[13][13] ), .ip2(n17378), .s(n17670), .op(n15608) );
  mux2_1 U19335 ( .ip1(\x[13][12] ), .ip2(n17379), .s(n17670), .op(n15607) );
  mux2_1 U19336 ( .ip1(\x[13][11] ), .ip2(n17380), .s(n17670), .op(n15606) );
  mux2_1 U19337 ( .ip1(\x[13][10] ), .ip2(n17381), .s(n17670), .op(n15605) );
  buf_1 U19338 ( .ip(n17670), .op(n17669) );
  mux2_1 U19339 ( .ip1(\x[13][9] ), .ip2(n17382), .s(n17669), .op(n15604) );
  mux2_1 U19340 ( .ip1(\x[13][8] ), .ip2(n17383), .s(n17670), .op(n15603) );
  mux2_1 U19341 ( .ip1(\x[13][7] ), .ip2(n17384), .s(n17669), .op(n15602) );
  mux2_1 U19342 ( .ip1(\x[13][6] ), .ip2(n17385), .s(n17670), .op(n15601) );
  mux2_1 U19343 ( .ip1(\x[13][5] ), .ip2(n17386), .s(n17669), .op(n15600) );
  mux2_1 U19344 ( .ip1(\x[13][4] ), .ip2(n17387), .s(n17670), .op(n15599) );
  mux2_1 U19345 ( .ip1(\x[13][3] ), .ip2(n17388), .s(n17669), .op(n15598) );
  mux2_1 U19346 ( .ip1(\x[13][2] ), .ip2(n17389), .s(n17669), .op(n15597) );
  mux2_1 U19347 ( .ip1(\x[13][1] ), .ip2(n17390), .s(n17669), .op(n15596) );
  mux2_1 U19348 ( .ip1(\x[13][0] ), .ip2(n17391), .s(n17669), .op(n15595) );
  buf_1 U19349 ( .ip(d[15]), .op(n17451) );
  nor2_1 U19350 ( .ip1(n17392), .ip2(n17404), .op(n17672) );
  mux2_1 U19351 ( .ip1(\x[12][15] ), .ip2(n17451), .s(n17672), .op(n15594) );
  buf_1 U19352 ( .ip(d[14]), .op(n17452) );
  mux2_1 U19353 ( .ip1(\x[12][14] ), .ip2(n17452), .s(n17672), .op(n15593) );
  buf_1 U19354 ( .ip(d[13]), .op(n17453) );
  mux2_1 U19355 ( .ip1(\x[12][13] ), .ip2(n17453), .s(n17672), .op(n15592) );
  buf_1 U19356 ( .ip(d[12]), .op(n17454) );
  mux2_1 U19357 ( .ip1(\x[12][12] ), .ip2(n17454), .s(n17672), .op(n15591) );
  buf_1 U19358 ( .ip(d[11]), .op(n17455) );
  mux2_1 U19359 ( .ip1(\x[12][11] ), .ip2(n17455), .s(n17672), .op(n15590) );
  buf_1 U19360 ( .ip(d[10]), .op(n17456) );
  mux2_1 U19361 ( .ip1(\x[12][10] ), .ip2(n17456), .s(n17672), .op(n15589) );
  buf_1 U19362 ( .ip(d[9]), .op(n17457) );
  buf_1 U19363 ( .ip(n17672), .op(n17671) );
  mux2_1 U19364 ( .ip1(\x[12][9] ), .ip2(n17457), .s(n17671), .op(n15588) );
  buf_1 U19365 ( .ip(d[8]), .op(n17458) );
  mux2_1 U19366 ( .ip1(\x[12][8] ), .ip2(n17458), .s(n17672), .op(n15587) );
  buf_1 U19367 ( .ip(d[7]), .op(n17459) );
  mux2_1 U19368 ( .ip1(\x[12][7] ), .ip2(n17459), .s(n17671), .op(n15586) );
  buf_1 U19369 ( .ip(d[6]), .op(n17461) );
  mux2_1 U19370 ( .ip1(\x[12][6] ), .ip2(n17461), .s(n17672), .op(n15585) );
  buf_1 U19371 ( .ip(d[5]), .op(n17462) );
  mux2_1 U19372 ( .ip1(\x[12][5] ), .ip2(n17462), .s(n17671), .op(n15584) );
  buf_1 U19373 ( .ip(d[4]), .op(n17463) );
  mux2_1 U19374 ( .ip1(\x[12][4] ), .ip2(n17463), .s(n17672), .op(n15583) );
  buf_1 U19375 ( .ip(d[3]), .op(n17464) );
  mux2_1 U19376 ( .ip1(\x[12][3] ), .ip2(n17464), .s(n17671), .op(n15582) );
  buf_1 U19377 ( .ip(d[2]), .op(n17465) );
  mux2_1 U19378 ( .ip1(\x[12][2] ), .ip2(n17465), .s(n17671), .op(n15581) );
  buf_1 U19379 ( .ip(d[1]), .op(n17466) );
  mux2_1 U19380 ( .ip1(\x[12][1] ), .ip2(n17466), .s(n17671), .op(n15580) );
  buf_1 U19381 ( .ip(d[0]), .op(n17468) );
  mux2_1 U19382 ( .ip1(\x[12][0] ), .ip2(n17468), .s(n17671), .op(n15579) );
  nor2_1 U19383 ( .ip1(n17393), .ip2(n17404), .op(n17674) );
  mux2_1 U19384 ( .ip1(\x[11][15] ), .ip2(n17451), .s(n17674), .op(n15578) );
  mux2_1 U19385 ( .ip1(\x[11][14] ), .ip2(n17452), .s(n17674), .op(n15577) );
  mux2_1 U19386 ( .ip1(\x[11][13] ), .ip2(n17453), .s(n17674), .op(n15576) );
  mux2_1 U19387 ( .ip1(\x[11][12] ), .ip2(n17454), .s(n17674), .op(n15575) );
  mux2_1 U19388 ( .ip1(\x[11][11] ), .ip2(n17455), .s(n17674), .op(n15574) );
  mux2_1 U19389 ( .ip1(\x[11][10] ), .ip2(n17456), .s(n17674), .op(n15573) );
  buf_1 U19390 ( .ip(n17674), .op(n17673) );
  mux2_1 U19391 ( .ip1(\x[11][9] ), .ip2(n17457), .s(n17673), .op(n15572) );
  mux2_1 U19392 ( .ip1(\x[11][8] ), .ip2(n17458), .s(n17674), .op(n15571) );
  mux2_1 U19393 ( .ip1(\x[11][7] ), .ip2(n17459), .s(n17673), .op(n15570) );
  mux2_1 U19394 ( .ip1(\x[11][6] ), .ip2(n17461), .s(n17674), .op(n15569) );
  mux2_1 U19395 ( .ip1(\x[11][5] ), .ip2(n17462), .s(n17673), .op(n15568) );
  mux2_1 U19396 ( .ip1(\x[11][4] ), .ip2(n17463), .s(n17674), .op(n15567) );
  mux2_1 U19397 ( .ip1(\x[11][3] ), .ip2(n17464), .s(n17673), .op(n15566) );
  mux2_1 U19398 ( .ip1(\x[11][2] ), .ip2(n17465), .s(n17673), .op(n15565) );
  mux2_1 U19399 ( .ip1(\x[11][1] ), .ip2(n17466), .s(n17673), .op(n15564) );
  mux2_1 U19400 ( .ip1(\x[11][0] ), .ip2(n17468), .s(n17673), .op(n15563) );
  nor2_1 U19401 ( .ip1(n17394), .ip2(n17404), .op(n17676) );
  mux2_1 U19402 ( .ip1(\x[10][15] ), .ip2(n17451), .s(n17676), .op(n15562) );
  mux2_1 U19403 ( .ip1(\x[10][14] ), .ip2(n17452), .s(n17676), .op(n15561) );
  mux2_1 U19404 ( .ip1(\x[10][13] ), .ip2(n17453), .s(n17676), .op(n15560) );
  mux2_1 U19405 ( .ip1(\x[10][12] ), .ip2(n17454), .s(n17676), .op(n15559) );
  mux2_1 U19406 ( .ip1(\x[10][11] ), .ip2(n17455), .s(n17676), .op(n15558) );
  mux2_1 U19407 ( .ip1(\x[10][10] ), .ip2(n17456), .s(n17676), .op(n15557) );
  buf_1 U19408 ( .ip(n17676), .op(n17675) );
  mux2_1 U19409 ( .ip1(\x[10][9] ), .ip2(n17457), .s(n17675), .op(n15556) );
  mux2_1 U19410 ( .ip1(\x[10][8] ), .ip2(n17458), .s(n17676), .op(n15555) );
  mux2_1 U19411 ( .ip1(\x[10][7] ), .ip2(n17459), .s(n17675), .op(n15554) );
  mux2_1 U19412 ( .ip1(\x[10][6] ), .ip2(n17461), .s(n17676), .op(n15553) );
  mux2_1 U19413 ( .ip1(\x[10][5] ), .ip2(n17462), .s(n17675), .op(n15552) );
  mux2_1 U19414 ( .ip1(\x[10][4] ), .ip2(n17463), .s(n17676), .op(n15551) );
  mux2_1 U19415 ( .ip1(\x[10][3] ), .ip2(n17464), .s(n17675), .op(n15550) );
  mux2_1 U19416 ( .ip1(\x[10][2] ), .ip2(n17465), .s(n17675), .op(n15549) );
  mux2_1 U19417 ( .ip1(\x[10][1] ), .ip2(n17466), .s(n17675), .op(n15548) );
  mux2_1 U19418 ( .ip1(\x[10][0] ), .ip2(n17468), .s(n17675), .op(n15547) );
  nor2_1 U19419 ( .ip1(n17395), .ip2(n17404), .op(n17678) );
  mux2_1 U19420 ( .ip1(\x[9][15] ), .ip2(n17451), .s(n17678), .op(n15546) );
  mux2_1 U19421 ( .ip1(\x[9][14] ), .ip2(n17452), .s(n17678), .op(n15545) );
  mux2_1 U19422 ( .ip1(\x[9][13] ), .ip2(n17453), .s(n17678), .op(n15544) );
  mux2_1 U19423 ( .ip1(\x[9][12] ), .ip2(n17454), .s(n17678), .op(n15543) );
  mux2_1 U19424 ( .ip1(\x[9][11] ), .ip2(n17455), .s(n17678), .op(n15542) );
  mux2_1 U19425 ( .ip1(\x[9][10] ), .ip2(n17456), .s(n17678), .op(n15541) );
  buf_1 U19426 ( .ip(n17678), .op(n17677) );
  mux2_1 U19427 ( .ip1(\x[9][9] ), .ip2(n17457), .s(n17677), .op(n15540) );
  mux2_1 U19428 ( .ip1(\x[9][8] ), .ip2(n17458), .s(n17678), .op(n15539) );
  mux2_1 U19429 ( .ip1(\x[9][7] ), .ip2(n17459), .s(n17677), .op(n15538) );
  mux2_1 U19430 ( .ip1(\x[9][6] ), .ip2(n17461), .s(n17678), .op(n15537) );
  mux2_1 U19431 ( .ip1(\x[9][5] ), .ip2(n17462), .s(n17677), .op(n15536) );
  mux2_1 U19432 ( .ip1(\x[9][4] ), .ip2(n17463), .s(n17678), .op(n15535) );
  mux2_1 U19433 ( .ip1(\x[9][3] ), .ip2(n17464), .s(n17677), .op(n15534) );
  mux2_1 U19434 ( .ip1(\x[9][2] ), .ip2(n17465), .s(n17677), .op(n15533) );
  mux2_1 U19435 ( .ip1(\x[9][1] ), .ip2(n17466), .s(n17677), .op(n15532) );
  mux2_1 U19436 ( .ip1(\x[9][0] ), .ip2(n17468), .s(n17677), .op(n15531) );
  nor2_1 U19437 ( .ip1(n17396), .ip2(n17404), .op(n17680) );
  mux2_1 U19438 ( .ip1(\x[8][15] ), .ip2(n17451), .s(n17680), .op(n15530) );
  mux2_1 U19439 ( .ip1(\x[8][14] ), .ip2(n17452), .s(n17680), .op(n15529) );
  mux2_1 U19440 ( .ip1(\x[8][13] ), .ip2(n17453), .s(n17680), .op(n15528) );
  mux2_1 U19441 ( .ip1(\x[8][12] ), .ip2(n17454), .s(n17680), .op(n15527) );
  mux2_1 U19442 ( .ip1(\x[8][11] ), .ip2(n17455), .s(n17680), .op(n15526) );
  mux2_1 U19443 ( .ip1(\x[8][10] ), .ip2(n17456), .s(n17680), .op(n15525) );
  buf_1 U19444 ( .ip(n17680), .op(n17679) );
  mux2_1 U19445 ( .ip1(\x[8][9] ), .ip2(n17457), .s(n17679), .op(n15524) );
  mux2_1 U19446 ( .ip1(\x[8][8] ), .ip2(n17458), .s(n17680), .op(n15523) );
  mux2_1 U19447 ( .ip1(\x[8][7] ), .ip2(n17459), .s(n17679), .op(n15522) );
  mux2_1 U19448 ( .ip1(\x[8][6] ), .ip2(n17461), .s(n17680), .op(n15521) );
  mux2_1 U19449 ( .ip1(\x[8][5] ), .ip2(n17462), .s(n17679), .op(n15520) );
  mux2_1 U19450 ( .ip1(\x[8][4] ), .ip2(n17463), .s(n17680), .op(n15519) );
  mux2_1 U19451 ( .ip1(\x[8][3] ), .ip2(n17464), .s(n17679), .op(n15518) );
  mux2_1 U19452 ( .ip1(\x[8][2] ), .ip2(n17465), .s(n17679), .op(n15517) );
  mux2_1 U19453 ( .ip1(\x[8][1] ), .ip2(n17466), .s(n17679), .op(n15516) );
  mux2_1 U19454 ( .ip1(\x[8][0] ), .ip2(n17468), .s(n17679), .op(n15515) );
  nor2_1 U19455 ( .ip1(n17397), .ip2(n17404), .op(n17682) );
  mux2_1 U19456 ( .ip1(\x[7][15] ), .ip2(n17451), .s(n17682), .op(n15514) );
  mux2_1 U19457 ( .ip1(\x[7][14] ), .ip2(n17452), .s(n17682), .op(n15513) );
  mux2_1 U19458 ( .ip1(\x[7][13] ), .ip2(n17453), .s(n17682), .op(n15512) );
  mux2_1 U19459 ( .ip1(\x[7][12] ), .ip2(n17454), .s(n17682), .op(n15511) );
  mux2_1 U19460 ( .ip1(\x[7][11] ), .ip2(n17455), .s(n17682), .op(n15510) );
  mux2_1 U19461 ( .ip1(\x[7][10] ), .ip2(n17456), .s(n17682), .op(n15509) );
  buf_1 U19462 ( .ip(n17682), .op(n17681) );
  mux2_1 U19463 ( .ip1(\x[7][9] ), .ip2(n17457), .s(n17681), .op(n15508) );
  mux2_1 U19464 ( .ip1(\x[7][8] ), .ip2(n17458), .s(n17682), .op(n15507) );
  mux2_1 U19465 ( .ip1(\x[7][7] ), .ip2(n17459), .s(n17681), .op(n15506) );
  mux2_1 U19466 ( .ip1(\x[7][6] ), .ip2(n17461), .s(n17682), .op(n15505) );
  mux2_1 U19467 ( .ip1(\x[7][5] ), .ip2(n17462), .s(n17681), .op(n15504) );
  mux2_1 U19468 ( .ip1(\x[7][4] ), .ip2(n17463), .s(n17682), .op(n15503) );
  mux2_1 U19469 ( .ip1(\x[7][3] ), .ip2(n17464), .s(n17681), .op(n15502) );
  mux2_1 U19470 ( .ip1(\x[7][2] ), .ip2(n17465), .s(n17681), .op(n15501) );
  mux2_1 U19471 ( .ip1(\x[7][1] ), .ip2(n17466), .s(n17681), .op(n15500) );
  mux2_1 U19472 ( .ip1(\x[7][0] ), .ip2(n17468), .s(n17681), .op(n15499) );
  nor2_1 U19473 ( .ip1(n17398), .ip2(n17404), .op(n17684) );
  mux2_1 U19474 ( .ip1(\x[6][15] ), .ip2(n17451), .s(n17684), .op(n15498) );
  mux2_1 U19475 ( .ip1(\x[6][14] ), .ip2(n17452), .s(n17684), .op(n15497) );
  mux2_1 U19476 ( .ip1(\x[6][13] ), .ip2(n17453), .s(n17684), .op(n15496) );
  mux2_1 U19477 ( .ip1(\x[6][12] ), .ip2(n17454), .s(n17684), .op(n15495) );
  mux2_1 U19478 ( .ip1(\x[6][11] ), .ip2(n17455), .s(n17684), .op(n15494) );
  mux2_1 U19479 ( .ip1(\x[6][10] ), .ip2(n17456), .s(n17684), .op(n15493) );
  buf_1 U19480 ( .ip(n17684), .op(n17683) );
  mux2_1 U19481 ( .ip1(\x[6][9] ), .ip2(n17457), .s(n17683), .op(n15492) );
  mux2_1 U19482 ( .ip1(\x[6][8] ), .ip2(n17458), .s(n17684), .op(n15491) );
  mux2_1 U19483 ( .ip1(\x[6][7] ), .ip2(n17459), .s(n17683), .op(n15490) );
  mux2_1 U19484 ( .ip1(\x[6][6] ), .ip2(n17461), .s(n17684), .op(n15489) );
  mux2_1 U19485 ( .ip1(\x[6][5] ), .ip2(n17462), .s(n17683), .op(n15488) );
  mux2_1 U19486 ( .ip1(\x[6][4] ), .ip2(n17463), .s(n17684), .op(n15487) );
  mux2_1 U19487 ( .ip1(\x[6][3] ), .ip2(n17464), .s(n17683), .op(n15486) );
  mux2_1 U19488 ( .ip1(\x[6][2] ), .ip2(n17465), .s(n17683), .op(n15485) );
  mux2_1 U19489 ( .ip1(\x[6][1] ), .ip2(n17466), .s(n17683), .op(n15484) );
  mux2_1 U19490 ( .ip1(\x[6][0] ), .ip2(n17468), .s(n17683), .op(n15483) );
  nor2_1 U19491 ( .ip1(n17399), .ip2(n17404), .op(n17686) );
  mux2_1 U19492 ( .ip1(\x[5][15] ), .ip2(n17451), .s(n17686), .op(n15482) );
  mux2_1 U19493 ( .ip1(\x[5][14] ), .ip2(n17452), .s(n17686), .op(n15481) );
  mux2_1 U19494 ( .ip1(\x[5][13] ), .ip2(n17453), .s(n17686), .op(n15480) );
  mux2_1 U19495 ( .ip1(\x[5][12] ), .ip2(n17454), .s(n17686), .op(n15479) );
  mux2_1 U19496 ( .ip1(\x[5][11] ), .ip2(n17455), .s(n17686), .op(n15478) );
  mux2_1 U19497 ( .ip1(\x[5][10] ), .ip2(n17456), .s(n17686), .op(n15477) );
  buf_1 U19498 ( .ip(n17686), .op(n17685) );
  mux2_1 U19499 ( .ip1(\x[5][9] ), .ip2(n17457), .s(n17685), .op(n15476) );
  mux2_1 U19500 ( .ip1(\x[5][8] ), .ip2(n17458), .s(n17686), .op(n15475) );
  mux2_1 U19501 ( .ip1(\x[5][7] ), .ip2(n17459), .s(n17685), .op(n15474) );
  mux2_1 U19502 ( .ip1(\x[5][6] ), .ip2(n17461), .s(n17686), .op(n15473) );
  mux2_1 U19503 ( .ip1(\x[5][5] ), .ip2(n17462), .s(n17685), .op(n15472) );
  mux2_1 U19504 ( .ip1(\x[5][4] ), .ip2(n17463), .s(n17686), .op(n15471) );
  mux2_1 U19505 ( .ip1(\x[5][3] ), .ip2(n17464), .s(n17685), .op(n15470) );
  mux2_1 U19506 ( .ip1(\x[5][2] ), .ip2(n17465), .s(n17685), .op(n15469) );
  mux2_1 U19507 ( .ip1(\x[5][1] ), .ip2(n17466), .s(n17685), .op(n15468) );
  mux2_1 U19508 ( .ip1(\x[5][0] ), .ip2(n17468), .s(n17685), .op(n15467) );
  nor2_1 U19509 ( .ip1(n17400), .ip2(n17404), .op(n17688) );
  mux2_1 U19510 ( .ip1(\x[4][15] ), .ip2(n17451), .s(n17688), .op(n15466) );
  mux2_1 U19511 ( .ip1(\x[4][14] ), .ip2(n17452), .s(n17688), .op(n15465) );
  mux2_1 U19512 ( .ip1(\x[4][13] ), .ip2(n17453), .s(n17688), .op(n15464) );
  mux2_1 U19513 ( .ip1(\x[4][12] ), .ip2(n17454), .s(n17688), .op(n15463) );
  mux2_1 U19514 ( .ip1(\x[4][11] ), .ip2(n17455), .s(n17688), .op(n15462) );
  mux2_1 U19515 ( .ip1(\x[4][10] ), .ip2(n17456), .s(n17688), .op(n15461) );
  buf_1 U19516 ( .ip(n17688), .op(n17687) );
  mux2_1 U19517 ( .ip1(\x[4][9] ), .ip2(n17457), .s(n17687), .op(n15460) );
  mux2_1 U19518 ( .ip1(\x[4][8] ), .ip2(n17458), .s(n17688), .op(n15459) );
  mux2_1 U19519 ( .ip1(\x[4][7] ), .ip2(n17459), .s(n17687), .op(n15458) );
  mux2_1 U19520 ( .ip1(\x[4][6] ), .ip2(n17461), .s(n17688), .op(n15457) );
  mux2_1 U19521 ( .ip1(\x[4][5] ), .ip2(n17462), .s(n17687), .op(n15456) );
  mux2_1 U19522 ( .ip1(\x[4][4] ), .ip2(n17463), .s(n17688), .op(n15455) );
  mux2_1 U19523 ( .ip1(\x[4][3] ), .ip2(n17464), .s(n17687), .op(n15454) );
  mux2_1 U19524 ( .ip1(\x[4][2] ), .ip2(n17465), .s(n17687), .op(n15453) );
  mux2_1 U19525 ( .ip1(\x[4][1] ), .ip2(n17466), .s(n17687), .op(n15452) );
  mux2_1 U19526 ( .ip1(\x[4][0] ), .ip2(n17468), .s(n17687), .op(n15451) );
  nor2_1 U19527 ( .ip1(n17401), .ip2(n17404), .op(n17690) );
  mux2_1 U19528 ( .ip1(\x[3][15] ), .ip2(n17451), .s(n17690), .op(n15450) );
  mux2_1 U19529 ( .ip1(\x[3][14] ), .ip2(n17452), .s(n17690), .op(n15449) );
  mux2_1 U19530 ( .ip1(\x[3][13] ), .ip2(n17453), .s(n17690), .op(n15448) );
  mux2_1 U19531 ( .ip1(\x[3][12] ), .ip2(n17454), .s(n17690), .op(n15447) );
  mux2_1 U19532 ( .ip1(\x[3][11] ), .ip2(n17455), .s(n17690), .op(n15446) );
  mux2_1 U19533 ( .ip1(\x[3][10] ), .ip2(n17456), .s(n17690), .op(n15445) );
  buf_1 U19534 ( .ip(n17690), .op(n17689) );
  mux2_1 U19535 ( .ip1(\x[3][9] ), .ip2(n17457), .s(n17689), .op(n15444) );
  mux2_1 U19536 ( .ip1(\x[3][8] ), .ip2(n17458), .s(n17690), .op(n15443) );
  mux2_1 U19537 ( .ip1(\x[3][7] ), .ip2(n17459), .s(n17689), .op(n15442) );
  mux2_1 U19538 ( .ip1(\x[3][6] ), .ip2(n17461), .s(n17690), .op(n15441) );
  mux2_1 U19539 ( .ip1(\x[3][5] ), .ip2(n17462), .s(n17689), .op(n15440) );
  mux2_1 U19540 ( .ip1(\x[3][4] ), .ip2(n17463), .s(n17690), .op(n15439) );
  mux2_1 U19541 ( .ip1(\x[3][3] ), .ip2(n17464), .s(n17689), .op(n15438) );
  mux2_1 U19542 ( .ip1(\x[3][2] ), .ip2(n17465), .s(n17689), .op(n15437) );
  mux2_1 U19543 ( .ip1(\x[3][1] ), .ip2(n17466), .s(n17689), .op(n15436) );
  mux2_1 U19544 ( .ip1(\x[3][0] ), .ip2(n17468), .s(n17689), .op(n15435) );
  nor2_1 U19545 ( .ip1(n17402), .ip2(n17404), .op(n17692) );
  mux2_1 U19546 ( .ip1(\x[2][15] ), .ip2(n17451), .s(n17692), .op(n15434) );
  mux2_1 U19547 ( .ip1(\x[2][14] ), .ip2(n17452), .s(n17692), .op(n15433) );
  mux2_1 U19548 ( .ip1(\x[2][13] ), .ip2(n17453), .s(n17692), .op(n15432) );
  mux2_1 U19549 ( .ip1(\x[2][12] ), .ip2(n17454), .s(n17692), .op(n15431) );
  mux2_1 U19550 ( .ip1(\x[2][11] ), .ip2(n17455), .s(n17692), .op(n15430) );
  mux2_1 U19551 ( .ip1(\x[2][10] ), .ip2(n17456), .s(n17692), .op(n15429) );
  buf_1 U19552 ( .ip(n17692), .op(n17691) );
  mux2_1 U19553 ( .ip1(\x[2][9] ), .ip2(n17457), .s(n17691), .op(n15428) );
  mux2_1 U19554 ( .ip1(\x[2][8] ), .ip2(n17458), .s(n17692), .op(n15427) );
  mux2_1 U19555 ( .ip1(\x[2][7] ), .ip2(n17459), .s(n17691), .op(n15426) );
  mux2_1 U19556 ( .ip1(\x[2][6] ), .ip2(n17461), .s(n17692), .op(n15425) );
  mux2_1 U19557 ( .ip1(\x[2][5] ), .ip2(n17462), .s(n17691), .op(n15424) );
  mux2_1 U19558 ( .ip1(\x[2][4] ), .ip2(n17463), .s(n17692), .op(n15423) );
  mux2_1 U19559 ( .ip1(\x[2][3] ), .ip2(n17464), .s(n17691), .op(n15422) );
  mux2_1 U19560 ( .ip1(\x[2][2] ), .ip2(n17465), .s(n17691), .op(n15421) );
  mux2_1 U19561 ( .ip1(\x[2][1] ), .ip2(n17466), .s(n17691), .op(n15420) );
  mux2_1 U19562 ( .ip1(\x[2][0] ), .ip2(n17468), .s(n17691), .op(n15419) );
  nor2_1 U19563 ( .ip1(n17403), .ip2(n17404), .op(n17694) );
  mux2_1 U19564 ( .ip1(\x[1][15] ), .ip2(n17451), .s(n17694), .op(n15418) );
  mux2_1 U19565 ( .ip1(\x[1][14] ), .ip2(n17452), .s(n17694), .op(n15417) );
  mux2_1 U19566 ( .ip1(\x[1][13] ), .ip2(n17453), .s(n17694), .op(n15416) );
  mux2_1 U19567 ( .ip1(\x[1][12] ), .ip2(n17454), .s(n17694), .op(n15415) );
  mux2_1 U19568 ( .ip1(\x[1][11] ), .ip2(n17455), .s(n17694), .op(n15414) );
  mux2_1 U19569 ( .ip1(\x[1][10] ), .ip2(n17456), .s(n17694), .op(n15413) );
  buf_1 U19570 ( .ip(n17694), .op(n17693) );
  mux2_1 U19571 ( .ip1(\x[1][9] ), .ip2(n17457), .s(n17693), .op(n15412) );
  mux2_1 U19572 ( .ip1(\x[1][8] ), .ip2(n17458), .s(n17694), .op(n15411) );
  mux2_1 U19573 ( .ip1(\x[1][7] ), .ip2(n17459), .s(n17693), .op(n15410) );
  mux2_1 U19574 ( .ip1(\x[1][6] ), .ip2(n17461), .s(n17694), .op(n15409) );
  mux2_1 U19575 ( .ip1(\x[1][5] ), .ip2(n17462), .s(n17693), .op(n15408) );
  mux2_1 U19576 ( .ip1(\x[1][4] ), .ip2(n17463), .s(n17694), .op(n15407) );
  mux2_1 U19577 ( .ip1(\x[1][3] ), .ip2(n17464), .s(n17693), .op(n15406) );
  mux2_1 U19578 ( .ip1(\x[1][2] ), .ip2(n17465), .s(n17693), .op(n15405) );
  mux2_1 U19579 ( .ip1(\x[1][1] ), .ip2(n17466), .s(n17693), .op(n15404) );
  mux2_1 U19580 ( .ip1(\x[1][0] ), .ip2(n17468), .s(n17693), .op(n15403) );
  nor2_1 U19581 ( .ip1(n17405), .ip2(n17404), .op(n17696) );
  mux2_1 U19582 ( .ip1(\x[0][15] ), .ip2(n17451), .s(n17696), .op(n15402) );
  mux2_1 U19583 ( .ip1(\x[0][14] ), .ip2(n17452), .s(n17696), .op(n15401) );
  mux2_1 U19584 ( .ip1(\x[0][13] ), .ip2(n17453), .s(n17696), .op(n15400) );
  mux2_1 U19585 ( .ip1(\x[0][12] ), .ip2(n17454), .s(n17696), .op(n15399) );
  mux2_1 U19586 ( .ip1(\x[0][11] ), .ip2(n17455), .s(n17696), .op(n15398) );
  mux2_1 U19587 ( .ip1(\x[0][10] ), .ip2(n17456), .s(n17696), .op(n15397) );
  buf_1 U19588 ( .ip(n17696), .op(n17695) );
  mux2_1 U19589 ( .ip1(\x[0][9] ), .ip2(n17457), .s(n17695), .op(n15396) );
  mux2_1 U19590 ( .ip1(\x[0][8] ), .ip2(n17458), .s(n17696), .op(n15395) );
  mux2_1 U19591 ( .ip1(\x[0][7] ), .ip2(n17459), .s(n17695), .op(n15394) );
  mux2_1 U19592 ( .ip1(\x[0][6] ), .ip2(n17461), .s(n17696), .op(n15393) );
  mux2_1 U19593 ( .ip1(\x[0][5] ), .ip2(n17462), .s(n17695), .op(n15392) );
  mux2_1 U19594 ( .ip1(\x[0][4] ), .ip2(n17463), .s(n17696), .op(n15391) );
  mux2_1 U19595 ( .ip1(\x[0][3] ), .ip2(n17464), .s(n17695), .op(n15390) );
  mux2_1 U19596 ( .ip1(\x[0][2] ), .ip2(n17465), .s(n17695), .op(n15389) );
  mux2_1 U19597 ( .ip1(\x[0][1] ), .ip2(n17466), .s(n17695), .op(n15388) );
  mux2_1 U19598 ( .ip1(\x[0][0] ), .ip2(n17468), .s(n17695), .op(n15387) );
  inv_1 U19599 ( .ip(done), .op(n17406) );
  nor3_1 U19600 ( .ip1(reset), .ip2(we), .ip3(n17406), .op(n26295) );
  inv_1 U19601 ( .ip(n26295), .op(n17408) );
  nand2_1 U19602 ( .ip1(we), .ip2(sig_ready), .op(n17407) );
  nand2_1 U19603 ( .ip1(n17408), .ip2(n17407), .op(n15386) );
  mux2_1 U19604 ( .ip1(\LUT[119][15] ), .ip2(n17451), .s(n17409), .op(n15385)
         );
  mux2_1 U19605 ( .ip1(\LUT[119][14] ), .ip2(n17452), .s(n17409), .op(n15384)
         );
  mux2_1 U19606 ( .ip1(\LUT[119][13] ), .ip2(n17453), .s(n17409), .op(n15383)
         );
  mux2_1 U19607 ( .ip1(\LUT[119][12] ), .ip2(n17454), .s(n17409), .op(n15382)
         );
  mux2_1 U19608 ( .ip1(\LUT[119][11] ), .ip2(n17455), .s(n17409), .op(n15381)
         );
  mux2_1 U19609 ( .ip1(\LUT[119][10] ), .ip2(n17456), .s(n17409), .op(n15380)
         );
  mux2_1 U19610 ( .ip1(\LUT[119][9] ), .ip2(n17457), .s(n17409), .op(n15379)
         );
  mux2_1 U19611 ( .ip1(\LUT[119][8] ), .ip2(n17458), .s(n17409), .op(n15378)
         );
  mux2_1 U19612 ( .ip1(\LUT[119][7] ), .ip2(n17459), .s(n17409), .op(n15377)
         );
  mux2_1 U19613 ( .ip1(\LUT[119][6] ), .ip2(n17461), .s(n17409), .op(n15376)
         );
  mux2_1 U19614 ( .ip1(\LUT[119][5] ), .ip2(n17462), .s(n17410), .op(n15375)
         );
  mux2_1 U19615 ( .ip1(\LUT[119][4] ), .ip2(n17463), .s(n17410), .op(n15374)
         );
  mux2_1 U19616 ( .ip1(\LUT[119][3] ), .ip2(n17464), .s(n17410), .op(n15373)
         );
  mux2_1 U19617 ( .ip1(\LUT[119][2] ), .ip2(n17465), .s(n17410), .op(n15372)
         );
  mux2_1 U19618 ( .ip1(\LUT[119][1] ), .ip2(n17466), .s(n17410), .op(n15371)
         );
  mux2_1 U19619 ( .ip1(\LUT[119][0] ), .ip2(n17468), .s(n17410), .op(n15370)
         );
  mux2_1 U19620 ( .ip1(\LUT[118][15] ), .ip2(n17451), .s(n17411), .op(n15369)
         );
  mux2_1 U19621 ( .ip1(\LUT[118][14] ), .ip2(n17452), .s(n17411), .op(n15368)
         );
  mux2_1 U19622 ( .ip1(\LUT[118][13] ), .ip2(n17453), .s(n17411), .op(n15367)
         );
  mux2_1 U19623 ( .ip1(\LUT[118][12] ), .ip2(n17454), .s(n17411), .op(n15366)
         );
  mux2_1 U19624 ( .ip1(\LUT[118][11] ), .ip2(n17455), .s(n17411), .op(n15365)
         );
  mux2_1 U19625 ( .ip1(\LUT[118][10] ), .ip2(n17456), .s(n17411), .op(n15364)
         );
  mux2_1 U19626 ( .ip1(\LUT[118][9] ), .ip2(n17457), .s(n17411), .op(n15363)
         );
  mux2_1 U19627 ( .ip1(\LUT[118][8] ), .ip2(n17458), .s(n17411), .op(n15362)
         );
  mux2_1 U19628 ( .ip1(\LUT[118][7] ), .ip2(n17459), .s(n17411), .op(n15361)
         );
  mux2_1 U19629 ( .ip1(\LUT[118][6] ), .ip2(n17461), .s(n17411), .op(n15360)
         );
  mux2_1 U19630 ( .ip1(\LUT[118][5] ), .ip2(n17462), .s(n17412), .op(n15359)
         );
  mux2_1 U19631 ( .ip1(\LUT[118][4] ), .ip2(n17463), .s(n17412), .op(n15358)
         );
  mux2_1 U19632 ( .ip1(\LUT[118][3] ), .ip2(n17464), .s(n17412), .op(n15357)
         );
  mux2_1 U19633 ( .ip1(\LUT[118][2] ), .ip2(n17465), .s(n17412), .op(n15356)
         );
  mux2_1 U19634 ( .ip1(\LUT[118][1] ), .ip2(n17466), .s(n17412), .op(n15355)
         );
  mux2_1 U19635 ( .ip1(\LUT[118][0] ), .ip2(n17468), .s(n17412), .op(n15354)
         );
  mux2_1 U19636 ( .ip1(\LUT[117][15] ), .ip2(n17451), .s(n17413), .op(n15353)
         );
  mux2_1 U19637 ( .ip1(\LUT[117][14] ), .ip2(n17452), .s(n17413), .op(n15352)
         );
  mux2_1 U19638 ( .ip1(\LUT[117][13] ), .ip2(n17453), .s(n17413), .op(n15351)
         );
  mux2_1 U19639 ( .ip1(\LUT[117][12] ), .ip2(n17454), .s(n17413), .op(n15350)
         );
  mux2_1 U19640 ( .ip1(\LUT[117][11] ), .ip2(n17455), .s(n17413), .op(n15349)
         );
  mux2_1 U19641 ( .ip1(\LUT[117][10] ), .ip2(n17456), .s(n17413), .op(n15348)
         );
  mux2_1 U19642 ( .ip1(\LUT[117][9] ), .ip2(n17457), .s(n17413), .op(n15347)
         );
  mux2_1 U19643 ( .ip1(\LUT[117][8] ), .ip2(n17458), .s(n17413), .op(n15346)
         );
  mux2_1 U19644 ( .ip1(\LUT[117][7] ), .ip2(n17459), .s(n17413), .op(n15345)
         );
  mux2_1 U19645 ( .ip1(\LUT[117][6] ), .ip2(n17461), .s(n17413), .op(n15344)
         );
  mux2_1 U19646 ( .ip1(\LUT[117][5] ), .ip2(n17462), .s(n17414), .op(n15343)
         );
  mux2_1 U19647 ( .ip1(\LUT[117][4] ), .ip2(n17463), .s(n17414), .op(n15342)
         );
  mux2_1 U19648 ( .ip1(\LUT[117][3] ), .ip2(n17464), .s(n17414), .op(n15341)
         );
  mux2_1 U19649 ( .ip1(\LUT[117][2] ), .ip2(n17465), .s(n17414), .op(n15340)
         );
  mux2_1 U19650 ( .ip1(\LUT[117][1] ), .ip2(n17466), .s(n17414), .op(n15339)
         );
  mux2_1 U19651 ( .ip1(\LUT[117][0] ), .ip2(n17468), .s(n17414), .op(n15338)
         );
  mux2_1 U19652 ( .ip1(\LUT[116][15] ), .ip2(n17451), .s(n17415), .op(n15337)
         );
  mux2_1 U19653 ( .ip1(\LUT[116][14] ), .ip2(n17452), .s(n17415), .op(n15336)
         );
  mux2_1 U19654 ( .ip1(\LUT[116][13] ), .ip2(n17453), .s(n17415), .op(n15335)
         );
  mux2_1 U19655 ( .ip1(\LUT[116][12] ), .ip2(n17454), .s(n17415), .op(n15334)
         );
  mux2_1 U19656 ( .ip1(\LUT[116][11] ), .ip2(n17455), .s(n17415), .op(n15333)
         );
  mux2_1 U19657 ( .ip1(\LUT[116][10] ), .ip2(n17456), .s(n17415), .op(n15332)
         );
  mux2_1 U19658 ( .ip1(\LUT[116][9] ), .ip2(n17457), .s(n17415), .op(n15331)
         );
  mux2_1 U19659 ( .ip1(\LUT[116][8] ), .ip2(n17458), .s(n17415), .op(n15330)
         );
  mux2_1 U19660 ( .ip1(\LUT[116][7] ), .ip2(n17459), .s(n17415), .op(n15329)
         );
  mux2_1 U19661 ( .ip1(\LUT[116][6] ), .ip2(n17461), .s(n17415), .op(n15328)
         );
  mux2_1 U19662 ( .ip1(\LUT[116][5] ), .ip2(n17462), .s(n17416), .op(n15327)
         );
  mux2_1 U19663 ( .ip1(\LUT[116][4] ), .ip2(n17463), .s(n17416), .op(n15326)
         );
  mux2_1 U19664 ( .ip1(\LUT[116][3] ), .ip2(n17464), .s(n17416), .op(n15325)
         );
  mux2_1 U19665 ( .ip1(\LUT[116][2] ), .ip2(n17465), .s(n17416), .op(n15324)
         );
  mux2_1 U19666 ( .ip1(\LUT[116][1] ), .ip2(n17466), .s(n17416), .op(n15323)
         );
  mux2_1 U19667 ( .ip1(\LUT[116][0] ), .ip2(n17468), .s(n17416), .op(n15322)
         );
  mux2_1 U19668 ( .ip1(\LUT[115][15] ), .ip2(n17451), .s(n17417), .op(n15321)
         );
  mux2_1 U19669 ( .ip1(\LUT[115][14] ), .ip2(n17452), .s(n17417), .op(n15320)
         );
  mux2_1 U19670 ( .ip1(\LUT[115][13] ), .ip2(n17453), .s(n17417), .op(n15319)
         );
  mux2_1 U19671 ( .ip1(\LUT[115][12] ), .ip2(n17454), .s(n17417), .op(n15318)
         );
  mux2_1 U19672 ( .ip1(\LUT[115][11] ), .ip2(n17455), .s(n17417), .op(n15317)
         );
  mux2_1 U19673 ( .ip1(\LUT[115][10] ), .ip2(n17456), .s(n17417), .op(n15316)
         );
  mux2_1 U19674 ( .ip1(\LUT[115][9] ), .ip2(n17457), .s(n17417), .op(n15315)
         );
  mux2_1 U19675 ( .ip1(\LUT[115][8] ), .ip2(n17458), .s(n17417), .op(n15314)
         );
  mux2_1 U19676 ( .ip1(\LUT[115][7] ), .ip2(n17459), .s(n17417), .op(n15313)
         );
  mux2_1 U19677 ( .ip1(\LUT[115][6] ), .ip2(n17461), .s(n17417), .op(n15312)
         );
  mux2_1 U19678 ( .ip1(\LUT[115][5] ), .ip2(n17462), .s(n17418), .op(n15311)
         );
  mux2_1 U19679 ( .ip1(\LUT[115][4] ), .ip2(n17463), .s(n17418), .op(n15310)
         );
  mux2_1 U19680 ( .ip1(\LUT[115][3] ), .ip2(n17464), .s(n17418), .op(n15309)
         );
  mux2_1 U19681 ( .ip1(\LUT[115][2] ), .ip2(n17465), .s(n17418), .op(n15308)
         );
  mux2_1 U19682 ( .ip1(\LUT[115][1] ), .ip2(n17466), .s(n17418), .op(n15307)
         );
  mux2_1 U19683 ( .ip1(\LUT[115][0] ), .ip2(n17468), .s(n17418), .op(n15306)
         );
  mux2_1 U19684 ( .ip1(\LUT[114][15] ), .ip2(n17451), .s(n17419), .op(n15305)
         );
  mux2_1 U19685 ( .ip1(\LUT[114][14] ), .ip2(n17452), .s(n17419), .op(n15304)
         );
  mux2_1 U19686 ( .ip1(\LUT[114][13] ), .ip2(n17453), .s(n17419), .op(n15303)
         );
  mux2_1 U19687 ( .ip1(\LUT[114][12] ), .ip2(n17454), .s(n17419), .op(n15302)
         );
  mux2_1 U19688 ( .ip1(\LUT[114][11] ), .ip2(n17455), .s(n17419), .op(n15301)
         );
  mux2_1 U19689 ( .ip1(\LUT[114][10] ), .ip2(n17456), .s(n17419), .op(n15300)
         );
  mux2_1 U19690 ( .ip1(\LUT[114][9] ), .ip2(n17457), .s(n17419), .op(n15299)
         );
  mux2_1 U19691 ( .ip1(\LUT[114][8] ), .ip2(n17458), .s(n17419), .op(n15298)
         );
  mux2_1 U19692 ( .ip1(\LUT[114][7] ), .ip2(n17459), .s(n17419), .op(n15297)
         );
  mux2_1 U19693 ( .ip1(\LUT[114][6] ), .ip2(n17461), .s(n17419), .op(n15296)
         );
  mux2_1 U19694 ( .ip1(\LUT[114][5] ), .ip2(n17462), .s(n17420), .op(n15295)
         );
  mux2_1 U19695 ( .ip1(\LUT[114][4] ), .ip2(n17463), .s(n17420), .op(n15294)
         );
  mux2_1 U19696 ( .ip1(\LUT[114][3] ), .ip2(n17464), .s(n17420), .op(n15293)
         );
  mux2_1 U19697 ( .ip1(\LUT[114][2] ), .ip2(n17465), .s(n17420), .op(n15292)
         );
  mux2_1 U19698 ( .ip1(\LUT[114][1] ), .ip2(n17466), .s(n17420), .op(n15291)
         );
  mux2_1 U19699 ( .ip1(\LUT[114][0] ), .ip2(n17468), .s(n17420), .op(n15290)
         );
  mux2_1 U19700 ( .ip1(\LUT[113][15] ), .ip2(n17451), .s(n17421), .op(n15289)
         );
  mux2_1 U19701 ( .ip1(\LUT[113][14] ), .ip2(n17452), .s(n17421), .op(n15288)
         );
  mux2_1 U19702 ( .ip1(\LUT[113][13] ), .ip2(n17453), .s(n17421), .op(n15287)
         );
  mux2_1 U19703 ( .ip1(\LUT[113][12] ), .ip2(n17454), .s(n17421), .op(n15286)
         );
  mux2_1 U19704 ( .ip1(\LUT[113][11] ), .ip2(n17455), .s(n17421), .op(n15285)
         );
  mux2_1 U19705 ( .ip1(\LUT[113][10] ), .ip2(n17456), .s(n17421), .op(n15284)
         );
  mux2_1 U19706 ( .ip1(\LUT[113][9] ), .ip2(n17457), .s(n17421), .op(n15283)
         );
  mux2_1 U19707 ( .ip1(\LUT[113][8] ), .ip2(n17458), .s(n17421), .op(n15282)
         );
  mux2_1 U19708 ( .ip1(\LUT[113][7] ), .ip2(n17459), .s(n17421), .op(n15281)
         );
  mux2_1 U19709 ( .ip1(\LUT[113][6] ), .ip2(n17461), .s(n17421), .op(n15280)
         );
  mux2_1 U19710 ( .ip1(\LUT[113][5] ), .ip2(n17462), .s(n17422), .op(n15279)
         );
  mux2_1 U19711 ( .ip1(\LUT[113][4] ), .ip2(n17463), .s(n17422), .op(n15278)
         );
  mux2_1 U19712 ( .ip1(\LUT[113][3] ), .ip2(n17464), .s(n17422), .op(n15277)
         );
  mux2_1 U19713 ( .ip1(\LUT[113][2] ), .ip2(n17465), .s(n17422), .op(n15276)
         );
  mux2_1 U19714 ( .ip1(\LUT[113][1] ), .ip2(n17466), .s(n17422), .op(n15275)
         );
  mux2_1 U19715 ( .ip1(\LUT[113][0] ), .ip2(n17468), .s(n17422), .op(n15274)
         );
  mux2_1 U19716 ( .ip1(\LUT[112][15] ), .ip2(n17451), .s(n17423), .op(n15273)
         );
  mux2_1 U19717 ( .ip1(\LUT[112][14] ), .ip2(n17452), .s(n17423), .op(n15272)
         );
  mux2_1 U19718 ( .ip1(\LUT[112][13] ), .ip2(n17453), .s(n17423), .op(n15271)
         );
  mux2_1 U19719 ( .ip1(\LUT[112][12] ), .ip2(n17454), .s(n17423), .op(n15270)
         );
  mux2_1 U19720 ( .ip1(\LUT[112][11] ), .ip2(n17455), .s(n17423), .op(n15269)
         );
  mux2_1 U19721 ( .ip1(\LUT[112][10] ), .ip2(n17456), .s(n17423), .op(n15268)
         );
  mux2_1 U19722 ( .ip1(\LUT[112][9] ), .ip2(n17457), .s(n17423), .op(n15267)
         );
  mux2_1 U19723 ( .ip1(\LUT[112][8] ), .ip2(n17458), .s(n17423), .op(n15266)
         );
  mux2_1 U19724 ( .ip1(\LUT[112][7] ), .ip2(n17459), .s(n17423), .op(n15265)
         );
  mux2_1 U19725 ( .ip1(\LUT[112][6] ), .ip2(n17461), .s(n17423), .op(n15264)
         );
  mux2_1 U19726 ( .ip1(\LUT[112][5] ), .ip2(n17462), .s(n17424), .op(n15263)
         );
  mux2_1 U19727 ( .ip1(\LUT[112][4] ), .ip2(n17463), .s(n17424), .op(n15262)
         );
  mux2_1 U19728 ( .ip1(\LUT[112][3] ), .ip2(n17464), .s(n17424), .op(n15261)
         );
  mux2_1 U19729 ( .ip1(\LUT[112][2] ), .ip2(n17465), .s(n17424), .op(n15260)
         );
  mux2_1 U19730 ( .ip1(\LUT[112][1] ), .ip2(n17466), .s(n17424), .op(n15259)
         );
  mux2_1 U19731 ( .ip1(\LUT[112][0] ), .ip2(n17468), .s(n17424), .op(n15258)
         );
  mux2_1 U19732 ( .ip1(\LUT[111][15] ), .ip2(n17451), .s(n17425), .op(n15257)
         );
  mux2_1 U19733 ( .ip1(\LUT[111][14] ), .ip2(n17452), .s(n17425), .op(n15256)
         );
  mux2_1 U19734 ( .ip1(\LUT[111][13] ), .ip2(n17453), .s(n17425), .op(n15255)
         );
  mux2_1 U19735 ( .ip1(\LUT[111][12] ), .ip2(n17454), .s(n17425), .op(n15254)
         );
  mux2_1 U19736 ( .ip1(\LUT[111][11] ), .ip2(n17455), .s(n17425), .op(n15253)
         );
  mux2_1 U19737 ( .ip1(\LUT[111][10] ), .ip2(n17456), .s(n17425), .op(n15252)
         );
  mux2_1 U19738 ( .ip1(\LUT[111][9] ), .ip2(n17457), .s(n17425), .op(n15251)
         );
  mux2_1 U19739 ( .ip1(\LUT[111][8] ), .ip2(n17458), .s(n17425), .op(n15250)
         );
  mux2_1 U19740 ( .ip1(\LUT[111][7] ), .ip2(n17459), .s(n17425), .op(n15249)
         );
  mux2_1 U19741 ( .ip1(\LUT[111][6] ), .ip2(n17461), .s(n17425), .op(n15248)
         );
  mux2_1 U19742 ( .ip1(\LUT[111][5] ), .ip2(n17462), .s(n17426), .op(n15247)
         );
  mux2_1 U19743 ( .ip1(\LUT[111][4] ), .ip2(n17463), .s(n17426), .op(n15246)
         );
  mux2_1 U19744 ( .ip1(\LUT[111][3] ), .ip2(n17464), .s(n17426), .op(n15245)
         );
  mux2_1 U19745 ( .ip1(\LUT[111][2] ), .ip2(n17465), .s(n17426), .op(n15244)
         );
  mux2_1 U19746 ( .ip1(\LUT[111][1] ), .ip2(n17466), .s(n17426), .op(n15243)
         );
  mux2_1 U19747 ( .ip1(\LUT[111][0] ), .ip2(n17468), .s(n17426), .op(n15242)
         );
  mux2_1 U19748 ( .ip1(\LUT[110][15] ), .ip2(n17451), .s(n17427), .op(n15241)
         );
  mux2_1 U19749 ( .ip1(\LUT[110][14] ), .ip2(n17452), .s(n17427), .op(n15240)
         );
  mux2_1 U19750 ( .ip1(\LUT[110][13] ), .ip2(n17453), .s(n17427), .op(n15239)
         );
  mux2_1 U19751 ( .ip1(\LUT[110][12] ), .ip2(n17454), .s(n17427), .op(n15238)
         );
  mux2_1 U19752 ( .ip1(\LUT[110][11] ), .ip2(n17455), .s(n17427), .op(n15237)
         );
  mux2_1 U19753 ( .ip1(\LUT[110][10] ), .ip2(n17456), .s(n17427), .op(n15236)
         );
  mux2_1 U19754 ( .ip1(\LUT[110][9] ), .ip2(n17457), .s(n17427), .op(n15235)
         );
  mux2_1 U19755 ( .ip1(\LUT[110][8] ), .ip2(n17458), .s(n17427), .op(n15234)
         );
  mux2_1 U19756 ( .ip1(\LUT[110][7] ), .ip2(n17459), .s(n17427), .op(n15233)
         );
  mux2_1 U19757 ( .ip1(\LUT[110][6] ), .ip2(n17461), .s(n17427), .op(n15232)
         );
  mux2_1 U19758 ( .ip1(\LUT[110][5] ), .ip2(n17462), .s(n17428), .op(n15231)
         );
  mux2_1 U19759 ( .ip1(\LUT[110][4] ), .ip2(n17463), .s(n17428), .op(n15230)
         );
  mux2_1 U19760 ( .ip1(\LUT[110][3] ), .ip2(n17464), .s(n17428), .op(n15229)
         );
  mux2_1 U19761 ( .ip1(\LUT[110][2] ), .ip2(n17465), .s(n17428), .op(n15228)
         );
  mux2_1 U19762 ( .ip1(\LUT[110][1] ), .ip2(n17466), .s(n17428), .op(n15227)
         );
  mux2_1 U19763 ( .ip1(\LUT[110][0] ), .ip2(n17468), .s(n17428), .op(n15226)
         );
  mux2_1 U19764 ( .ip1(\LUT[109][15] ), .ip2(n17451), .s(n17429), .op(n15225)
         );
  mux2_1 U19765 ( .ip1(\LUT[109][14] ), .ip2(n17452), .s(n17429), .op(n15224)
         );
  mux2_1 U19766 ( .ip1(\LUT[109][13] ), .ip2(n17453), .s(n17429), .op(n15223)
         );
  mux2_1 U19767 ( .ip1(\LUT[109][12] ), .ip2(n17454), .s(n17429), .op(n15222)
         );
  mux2_1 U19768 ( .ip1(\LUT[109][11] ), .ip2(n17455), .s(n17429), .op(n15221)
         );
  mux2_1 U19769 ( .ip1(\LUT[109][10] ), .ip2(n17456), .s(n17429), .op(n15220)
         );
  mux2_1 U19770 ( .ip1(\LUT[109][9] ), .ip2(n17457), .s(n17429), .op(n15219)
         );
  mux2_1 U19771 ( .ip1(\LUT[109][8] ), .ip2(n17458), .s(n17429), .op(n15218)
         );
  mux2_1 U19772 ( .ip1(\LUT[109][7] ), .ip2(n17459), .s(n17429), .op(n15217)
         );
  mux2_1 U19773 ( .ip1(\LUT[109][6] ), .ip2(n17461), .s(n17429), .op(n15216)
         );
  mux2_1 U19774 ( .ip1(\LUT[109][5] ), .ip2(n17462), .s(n17430), .op(n15215)
         );
  mux2_1 U19775 ( .ip1(\LUT[109][4] ), .ip2(n17463), .s(n17430), .op(n15214)
         );
  mux2_1 U19776 ( .ip1(\LUT[109][3] ), .ip2(n17464), .s(n17430), .op(n15213)
         );
  mux2_1 U19777 ( .ip1(\LUT[109][2] ), .ip2(n17465), .s(n17430), .op(n15212)
         );
  mux2_1 U19778 ( .ip1(\LUT[109][1] ), .ip2(n17466), .s(n17430), .op(n15211)
         );
  mux2_1 U19779 ( .ip1(\LUT[109][0] ), .ip2(n17468), .s(n17430), .op(n15210)
         );
  mux2_1 U19780 ( .ip1(\LUT[108][15] ), .ip2(n17451), .s(n17431), .op(n15209)
         );
  mux2_1 U19781 ( .ip1(\LUT[108][14] ), .ip2(n17452), .s(n17431), .op(n15208)
         );
  mux2_1 U19782 ( .ip1(\LUT[108][13] ), .ip2(n17453), .s(n17431), .op(n15207)
         );
  mux2_1 U19783 ( .ip1(\LUT[108][12] ), .ip2(n17454), .s(n17431), .op(n15206)
         );
  mux2_1 U19784 ( .ip1(\LUT[108][11] ), .ip2(n17455), .s(n17431), .op(n15205)
         );
  mux2_1 U19785 ( .ip1(\LUT[108][10] ), .ip2(n17456), .s(n17431), .op(n15204)
         );
  mux2_1 U19786 ( .ip1(\LUT[108][9] ), .ip2(n17457), .s(n17431), .op(n15203)
         );
  mux2_1 U19787 ( .ip1(\LUT[108][8] ), .ip2(n17458), .s(n17431), .op(n15202)
         );
  mux2_1 U19788 ( .ip1(\LUT[108][7] ), .ip2(n17459), .s(n17431), .op(n15201)
         );
  mux2_1 U19789 ( .ip1(\LUT[108][6] ), .ip2(n17461), .s(n17431), .op(n15200)
         );
  mux2_1 U19790 ( .ip1(\LUT[108][5] ), .ip2(n17462), .s(n17432), .op(n15199)
         );
  mux2_1 U19791 ( .ip1(\LUT[108][4] ), .ip2(n17463), .s(n17432), .op(n15198)
         );
  mux2_1 U19792 ( .ip1(\LUT[108][3] ), .ip2(n17464), .s(n17432), .op(n15197)
         );
  mux2_1 U19793 ( .ip1(\LUT[108][2] ), .ip2(n17465), .s(n17432), .op(n15196)
         );
  mux2_1 U19794 ( .ip1(\LUT[108][1] ), .ip2(n17466), .s(n17432), .op(n15195)
         );
  mux2_1 U19795 ( .ip1(\LUT[108][0] ), .ip2(n17468), .s(n17432), .op(n15194)
         );
  mux2_1 U19796 ( .ip1(\LUT[107][15] ), .ip2(n17451), .s(n17433), .op(n15193)
         );
  mux2_1 U19797 ( .ip1(\LUT[107][14] ), .ip2(n17452), .s(n17433), .op(n15192)
         );
  mux2_1 U19798 ( .ip1(\LUT[107][13] ), .ip2(n17453), .s(n17433), .op(n15191)
         );
  mux2_1 U19799 ( .ip1(\LUT[107][12] ), .ip2(n17454), .s(n17433), .op(n15190)
         );
  mux2_1 U19800 ( .ip1(\LUT[107][11] ), .ip2(n17455), .s(n17433), .op(n15189)
         );
  mux2_1 U19801 ( .ip1(\LUT[107][10] ), .ip2(n17456), .s(n17433), .op(n15188)
         );
  mux2_1 U19802 ( .ip1(\LUT[107][9] ), .ip2(n17457), .s(n17433), .op(n15187)
         );
  mux2_1 U19803 ( .ip1(\LUT[107][8] ), .ip2(n17458), .s(n17433), .op(n15186)
         );
  mux2_1 U19804 ( .ip1(\LUT[107][7] ), .ip2(n17459), .s(n17433), .op(n15185)
         );
  mux2_1 U19805 ( .ip1(\LUT[107][6] ), .ip2(n17461), .s(n17433), .op(n15184)
         );
  mux2_1 U19806 ( .ip1(\LUT[107][5] ), .ip2(n17462), .s(n17434), .op(n15183)
         );
  mux2_1 U19807 ( .ip1(\LUT[107][4] ), .ip2(n17463), .s(n17434), .op(n15182)
         );
  mux2_1 U19808 ( .ip1(\LUT[107][3] ), .ip2(n17464), .s(n17434), .op(n15181)
         );
  mux2_1 U19809 ( .ip1(\LUT[107][2] ), .ip2(n17465), .s(n17434), .op(n15180)
         );
  mux2_1 U19810 ( .ip1(\LUT[107][1] ), .ip2(n17466), .s(n17434), .op(n15179)
         );
  mux2_1 U19811 ( .ip1(\LUT[107][0] ), .ip2(n17468), .s(n17434), .op(n15178)
         );
  mux2_1 U19812 ( .ip1(\LUT[106][15] ), .ip2(n17451), .s(n17435), .op(n15177)
         );
  mux2_1 U19813 ( .ip1(\LUT[106][14] ), .ip2(n17452), .s(n17435), .op(n15176)
         );
  mux2_1 U19814 ( .ip1(\LUT[106][13] ), .ip2(n17453), .s(n17435), .op(n15175)
         );
  mux2_1 U19815 ( .ip1(\LUT[106][12] ), .ip2(n17454), .s(n17435), .op(n15174)
         );
  mux2_1 U19816 ( .ip1(\LUT[106][11] ), .ip2(n17455), .s(n17435), .op(n15173)
         );
  mux2_1 U19817 ( .ip1(\LUT[106][10] ), .ip2(n17456), .s(n17435), .op(n15172)
         );
  mux2_1 U19818 ( .ip1(\LUT[106][9] ), .ip2(n17457), .s(n17435), .op(n15171)
         );
  mux2_1 U19819 ( .ip1(\LUT[106][8] ), .ip2(n17458), .s(n17435), .op(n15170)
         );
  mux2_1 U19820 ( .ip1(\LUT[106][7] ), .ip2(n17459), .s(n17435), .op(n15169)
         );
  mux2_1 U19821 ( .ip1(\LUT[106][6] ), .ip2(n17461), .s(n17435), .op(n15168)
         );
  mux2_1 U19822 ( .ip1(\LUT[106][5] ), .ip2(n17462), .s(n17436), .op(n15167)
         );
  mux2_1 U19823 ( .ip1(\LUT[106][4] ), .ip2(n17463), .s(n17436), .op(n15166)
         );
  mux2_1 U19824 ( .ip1(\LUT[106][3] ), .ip2(n17464), .s(n17436), .op(n15165)
         );
  mux2_1 U19825 ( .ip1(\LUT[106][2] ), .ip2(n17465), .s(n17436), .op(n15164)
         );
  mux2_1 U19826 ( .ip1(\LUT[106][1] ), .ip2(n17466), .s(n17436), .op(n15163)
         );
  mux2_1 U19827 ( .ip1(\LUT[106][0] ), .ip2(n17468), .s(n17436), .op(n15162)
         );
  mux2_1 U19828 ( .ip1(\LUT[105][15] ), .ip2(n17451), .s(n17437), .op(n15161)
         );
  mux2_1 U19829 ( .ip1(\LUT[105][14] ), .ip2(n17452), .s(n17437), .op(n15160)
         );
  mux2_1 U19830 ( .ip1(\LUT[105][13] ), .ip2(n17453), .s(n17437), .op(n15159)
         );
  mux2_1 U19831 ( .ip1(\LUT[105][12] ), .ip2(n17454), .s(n17437), .op(n15158)
         );
  mux2_1 U19832 ( .ip1(\LUT[105][11] ), .ip2(n17455), .s(n17437), .op(n15157)
         );
  mux2_1 U19833 ( .ip1(\LUT[105][10] ), .ip2(n17456), .s(n17437), .op(n15156)
         );
  mux2_1 U19834 ( .ip1(\LUT[105][9] ), .ip2(n17457), .s(n17437), .op(n15155)
         );
  mux2_1 U19835 ( .ip1(\LUT[105][8] ), .ip2(n17458), .s(n17437), .op(n15154)
         );
  mux2_1 U19836 ( .ip1(\LUT[105][7] ), .ip2(n17459), .s(n17437), .op(n15153)
         );
  mux2_1 U19837 ( .ip1(\LUT[105][6] ), .ip2(n17461), .s(n17437), .op(n15152)
         );
  mux2_1 U19838 ( .ip1(\LUT[105][5] ), .ip2(n17462), .s(n17438), .op(n15151)
         );
  mux2_1 U19839 ( .ip1(\LUT[105][4] ), .ip2(n17463), .s(n17438), .op(n15150)
         );
  mux2_1 U19840 ( .ip1(\LUT[105][3] ), .ip2(n17464), .s(n17438), .op(n15149)
         );
  mux2_1 U19841 ( .ip1(\LUT[105][2] ), .ip2(n17465), .s(n17438), .op(n15148)
         );
  mux2_1 U19842 ( .ip1(\LUT[105][1] ), .ip2(n17466), .s(n17438), .op(n15147)
         );
  mux2_1 U19843 ( .ip1(\LUT[105][0] ), .ip2(n17468), .s(n17438), .op(n15146)
         );
  mux2_1 U19844 ( .ip1(\LUT[104][15] ), .ip2(n17451), .s(n17439), .op(n15145)
         );
  mux2_1 U19845 ( .ip1(\LUT[104][14] ), .ip2(n17452), .s(n17439), .op(n15144)
         );
  mux2_1 U19846 ( .ip1(\LUT[104][13] ), .ip2(n17453), .s(n17439), .op(n15143)
         );
  mux2_1 U19847 ( .ip1(\LUT[104][12] ), .ip2(n17454), .s(n17439), .op(n15142)
         );
  mux2_1 U19848 ( .ip1(\LUT[104][11] ), .ip2(n17455), .s(n17439), .op(n15141)
         );
  mux2_1 U19849 ( .ip1(\LUT[104][10] ), .ip2(n17456), .s(n17439), .op(n15140)
         );
  mux2_1 U19850 ( .ip1(\LUT[104][9] ), .ip2(n17457), .s(n17439), .op(n15139)
         );
  mux2_1 U19851 ( .ip1(\LUT[104][8] ), .ip2(n17458), .s(n17439), .op(n15138)
         );
  mux2_1 U19852 ( .ip1(\LUT[104][7] ), .ip2(n17459), .s(n17439), .op(n15137)
         );
  mux2_1 U19853 ( .ip1(\LUT[104][6] ), .ip2(n17461), .s(n17439), .op(n15136)
         );
  mux2_1 U19854 ( .ip1(\LUT[104][5] ), .ip2(n17462), .s(n17440), .op(n15135)
         );
  mux2_1 U19855 ( .ip1(\LUT[104][4] ), .ip2(n17463), .s(n17440), .op(n15134)
         );
  mux2_1 U19856 ( .ip1(\LUT[104][3] ), .ip2(n17464), .s(n17440), .op(n15133)
         );
  mux2_1 U19857 ( .ip1(\LUT[104][2] ), .ip2(n17465), .s(n17440), .op(n15132)
         );
  mux2_1 U19858 ( .ip1(\LUT[104][1] ), .ip2(n17466), .s(n17440), .op(n15131)
         );
  mux2_1 U19859 ( .ip1(\LUT[104][0] ), .ip2(n17468), .s(n17440), .op(n15130)
         );
  mux2_1 U19860 ( .ip1(\LUT[103][15] ), .ip2(n17451), .s(n17441), .op(n15129)
         );
  mux2_1 U19861 ( .ip1(\LUT[103][14] ), .ip2(n17452), .s(n17441), .op(n15128)
         );
  mux2_1 U19862 ( .ip1(\LUT[103][13] ), .ip2(n17453), .s(n17441), .op(n15127)
         );
  mux2_1 U19863 ( .ip1(\LUT[103][12] ), .ip2(n17454), .s(n17441), .op(n15126)
         );
  mux2_1 U19864 ( .ip1(\LUT[103][11] ), .ip2(n17455), .s(n17441), .op(n15125)
         );
  mux2_1 U19865 ( .ip1(\LUT[103][10] ), .ip2(n17456), .s(n17441), .op(n15124)
         );
  mux2_1 U19866 ( .ip1(\LUT[103][9] ), .ip2(n17457), .s(n17441), .op(n15123)
         );
  mux2_1 U19867 ( .ip1(\LUT[103][8] ), .ip2(n17458), .s(n17441), .op(n15122)
         );
  mux2_1 U19868 ( .ip1(\LUT[103][7] ), .ip2(n17459), .s(n17441), .op(n15121)
         );
  mux2_1 U19869 ( .ip1(\LUT[103][6] ), .ip2(n17461), .s(n17441), .op(n15120)
         );
  mux2_1 U19870 ( .ip1(\LUT[103][5] ), .ip2(n17462), .s(n17442), .op(n15119)
         );
  mux2_1 U19871 ( .ip1(\LUT[103][4] ), .ip2(n17463), .s(n17442), .op(n15118)
         );
  mux2_1 U19872 ( .ip1(\LUT[103][3] ), .ip2(n17464), .s(n17442), .op(n15117)
         );
  mux2_1 U19873 ( .ip1(\LUT[103][2] ), .ip2(n17465), .s(n17442), .op(n15116)
         );
  mux2_1 U19874 ( .ip1(\LUT[103][1] ), .ip2(n17466), .s(n17442), .op(n15115)
         );
  mux2_1 U19875 ( .ip1(\LUT[103][0] ), .ip2(n17468), .s(n17442), .op(n15114)
         );
  mux2_1 U19876 ( .ip1(\LUT[102][15] ), .ip2(n17451), .s(n17443), .op(n15113)
         );
  mux2_1 U19877 ( .ip1(\LUT[102][14] ), .ip2(n17452), .s(n17443), .op(n15112)
         );
  mux2_1 U19878 ( .ip1(\LUT[102][13] ), .ip2(n17453), .s(n17443), .op(n15111)
         );
  mux2_1 U19879 ( .ip1(\LUT[102][12] ), .ip2(n17454), .s(n17443), .op(n15110)
         );
  mux2_1 U19880 ( .ip1(\LUT[102][11] ), .ip2(n17455), .s(n17443), .op(n15109)
         );
  mux2_1 U19881 ( .ip1(\LUT[102][10] ), .ip2(n17456), .s(n17443), .op(n15108)
         );
  mux2_1 U19882 ( .ip1(\LUT[102][9] ), .ip2(n17457), .s(n17443), .op(n15107)
         );
  mux2_1 U19883 ( .ip1(\LUT[102][8] ), .ip2(n17458), .s(n17443), .op(n15106)
         );
  mux2_1 U19884 ( .ip1(\LUT[102][7] ), .ip2(n17459), .s(n17443), .op(n15105)
         );
  mux2_1 U19885 ( .ip1(\LUT[102][6] ), .ip2(n17461), .s(n17443), .op(n15104)
         );
  mux2_1 U19886 ( .ip1(\LUT[102][5] ), .ip2(n17462), .s(n17444), .op(n15103)
         );
  mux2_1 U19887 ( .ip1(\LUT[102][4] ), .ip2(n17463), .s(n17444), .op(n15102)
         );
  mux2_1 U19888 ( .ip1(\LUT[102][3] ), .ip2(n17464), .s(n17444), .op(n15101)
         );
  mux2_1 U19889 ( .ip1(\LUT[102][2] ), .ip2(n17465), .s(n17444), .op(n15100)
         );
  mux2_1 U19890 ( .ip1(\LUT[102][1] ), .ip2(n17466), .s(n17444), .op(n15099)
         );
  mux2_1 U19891 ( .ip1(\LUT[102][0] ), .ip2(n17468), .s(n17444), .op(n15098)
         );
  mux2_1 U19892 ( .ip1(\LUT[101][15] ), .ip2(d[15]), .s(n17445), .op(n15097)
         );
  mux2_1 U19893 ( .ip1(\LUT[101][14] ), .ip2(d[14]), .s(n17445), .op(n15096)
         );
  mux2_1 U19894 ( .ip1(\LUT[101][13] ), .ip2(d[13]), .s(n17445), .op(n15095)
         );
  mux2_1 U19895 ( .ip1(\LUT[101][12] ), .ip2(d[12]), .s(n17445), .op(n15094)
         );
  mux2_1 U19896 ( .ip1(\LUT[101][11] ), .ip2(d[11]), .s(n17445), .op(n15093)
         );
  mux2_1 U19897 ( .ip1(\LUT[101][10] ), .ip2(d[10]), .s(n17445), .op(n15092)
         );
  mux2_1 U19898 ( .ip1(\LUT[101][9] ), .ip2(d[9]), .s(n17445), .op(n15091) );
  mux2_1 U19899 ( .ip1(\LUT[101][8] ), .ip2(d[8]), .s(n17445), .op(n15090) );
  mux2_1 U19900 ( .ip1(\LUT[101][7] ), .ip2(d[7]), .s(n17445), .op(n15089) );
  mux2_1 U19901 ( .ip1(\LUT[101][6] ), .ip2(d[6]), .s(n17445), .op(n15088) );
  mux2_1 U19902 ( .ip1(\LUT[101][5] ), .ip2(d[5]), .s(n17446), .op(n15087) );
  mux2_1 U19903 ( .ip1(\LUT[101][4] ), .ip2(d[4]), .s(n17446), .op(n15086) );
  mux2_1 U19904 ( .ip1(\LUT[101][3] ), .ip2(d[3]), .s(n17446), .op(n15085) );
  mux2_1 U19905 ( .ip1(\LUT[101][2] ), .ip2(d[2]), .s(n17446), .op(n15084) );
  mux2_1 U19906 ( .ip1(\LUT[101][1] ), .ip2(d[1]), .s(n17446), .op(n15083) );
  mux2_1 U19907 ( .ip1(\LUT[101][0] ), .ip2(d[0]), .s(n17446), .op(n15082) );
  mux2_1 U19908 ( .ip1(\LUT[100][15] ), .ip2(n17451), .s(n17447), .op(n15081)
         );
  mux2_1 U19909 ( .ip1(\LUT[100][14] ), .ip2(n17452), .s(n17447), .op(n15080)
         );
  mux2_1 U19910 ( .ip1(\LUT[100][13] ), .ip2(n17453), .s(n17447), .op(n15079)
         );
  mux2_1 U19911 ( .ip1(\LUT[100][12] ), .ip2(n17454), .s(n17447), .op(n15078)
         );
  mux2_1 U19912 ( .ip1(\LUT[100][11] ), .ip2(n17455), .s(n17447), .op(n15077)
         );
  mux2_1 U19913 ( .ip1(\LUT[100][10] ), .ip2(n17456), .s(n17447), .op(n15076)
         );
  mux2_1 U19914 ( .ip1(\LUT[100][9] ), .ip2(n17457), .s(n17447), .op(n15075)
         );
  mux2_1 U19915 ( .ip1(\LUT[100][8] ), .ip2(n17458), .s(n17447), .op(n15074)
         );
  mux2_1 U19916 ( .ip1(\LUT[100][7] ), .ip2(n17459), .s(n17447), .op(n15073)
         );
  mux2_1 U19917 ( .ip1(\LUT[100][6] ), .ip2(n17461), .s(n17447), .op(n15072)
         );
  mux2_1 U19918 ( .ip1(\LUT[100][5] ), .ip2(n17462), .s(n17448), .op(n15071)
         );
  mux2_1 U19919 ( .ip1(\LUT[100][4] ), .ip2(n17463), .s(n17448), .op(n15070)
         );
  mux2_1 U19920 ( .ip1(\LUT[100][3] ), .ip2(n17464), .s(n17448), .op(n15069)
         );
  mux2_1 U19921 ( .ip1(\LUT[100][2] ), .ip2(n17465), .s(n17448), .op(n15068)
         );
  mux2_1 U19922 ( .ip1(\LUT[100][1] ), .ip2(n17466), .s(n17448), .op(n15067)
         );
  mux2_1 U19923 ( .ip1(\LUT[100][0] ), .ip2(n17468), .s(n17448), .op(n15066)
         );
  mux2_1 U19924 ( .ip1(\LUT[99][15] ), .ip2(d[15]), .s(n17449), .op(n15065) );
  mux2_1 U19925 ( .ip1(\LUT[99][14] ), .ip2(d[14]), .s(n17449), .op(n15064) );
  mux2_1 U19926 ( .ip1(\LUT[99][13] ), .ip2(d[13]), .s(n17449), .op(n15063) );
  mux2_1 U19927 ( .ip1(\LUT[99][12] ), .ip2(d[12]), .s(n17449), .op(n15062) );
  mux2_1 U19928 ( .ip1(\LUT[99][11] ), .ip2(d[11]), .s(n17449), .op(n15061) );
  mux2_1 U19929 ( .ip1(\LUT[99][10] ), .ip2(d[10]), .s(n17449), .op(n15060) );
  mux2_1 U19930 ( .ip1(\LUT[99][9] ), .ip2(d[9]), .s(n17449), .op(n15059) );
  mux2_1 U19931 ( .ip1(\LUT[99][8] ), .ip2(d[8]), .s(n17449), .op(n15058) );
  mux2_1 U19932 ( .ip1(\LUT[99][7] ), .ip2(d[7]), .s(n17449), .op(n15057) );
  mux2_1 U19933 ( .ip1(\LUT[99][6] ), .ip2(d[6]), .s(n17449), .op(n15056) );
  mux2_1 U19934 ( .ip1(\LUT[99][5] ), .ip2(d[5]), .s(n17450), .op(n15055) );
  mux2_1 U19935 ( .ip1(\LUT[99][4] ), .ip2(d[4]), .s(n17450), .op(n15054) );
  mux2_1 U19936 ( .ip1(\LUT[99][3] ), .ip2(d[3]), .s(n17450), .op(n15053) );
  mux2_1 U19937 ( .ip1(\LUT[99][2] ), .ip2(d[2]), .s(n17450), .op(n15052) );
  mux2_1 U19938 ( .ip1(\LUT[99][1] ), .ip2(d[1]), .s(n17450), .op(n15051) );
  mux2_1 U19939 ( .ip1(\LUT[99][0] ), .ip2(d[0]), .s(n17450), .op(n15050) );
  mux2_1 U19940 ( .ip1(\LUT[98][15] ), .ip2(n17451), .s(n17460), .op(n15049)
         );
  mux2_1 U19941 ( .ip1(\LUT[98][14] ), .ip2(n17452), .s(n17460), .op(n15048)
         );
  mux2_1 U19942 ( .ip1(\LUT[98][13] ), .ip2(n17453), .s(n17460), .op(n15047)
         );
  mux2_1 U19943 ( .ip1(\LUT[98][12] ), .ip2(n17454), .s(n17460), .op(n15046)
         );
  mux2_1 U19944 ( .ip1(\LUT[98][11] ), .ip2(n17455), .s(n17460), .op(n15045)
         );
  mux2_1 U19945 ( .ip1(\LUT[98][10] ), .ip2(n17456), .s(n17460), .op(n15044)
         );
  mux2_1 U19946 ( .ip1(\LUT[98][9] ), .ip2(n17457), .s(n17460), .op(n15043) );
  mux2_1 U19947 ( .ip1(\LUT[98][8] ), .ip2(n17458), .s(n17460), .op(n15042) );
  mux2_1 U19948 ( .ip1(\LUT[98][7] ), .ip2(n17459), .s(n17460), .op(n15041) );
  mux2_1 U19949 ( .ip1(\LUT[98][6] ), .ip2(n17461), .s(n17460), .op(n15040) );
  mux2_1 U19950 ( .ip1(\LUT[98][5] ), .ip2(n17462), .s(n17467), .op(n15039) );
  mux2_1 U19951 ( .ip1(\LUT[98][4] ), .ip2(n17463), .s(n17467), .op(n15038) );
  mux2_1 U19952 ( .ip1(\LUT[98][3] ), .ip2(n17464), .s(n17467), .op(n15037) );
  mux2_1 U19953 ( .ip1(\LUT[98][2] ), .ip2(n17465), .s(n17467), .op(n15036) );
  mux2_1 U19954 ( .ip1(\LUT[98][1] ), .ip2(n17466), .s(n17467), .op(n15035) );
  mux2_1 U19955 ( .ip1(\LUT[98][0] ), .ip2(n17468), .s(n17467), .op(n15034) );
  mux2_1 U19956 ( .ip1(\LUT[97][15] ), .ip2(d[15]), .s(n17469), .op(n15033) );
  mux2_1 U19957 ( .ip1(\LUT[97][14] ), .ip2(d[14]), .s(n17469), .op(n15032) );
  mux2_1 U19958 ( .ip1(\LUT[97][13] ), .ip2(d[13]), .s(n17469), .op(n15031) );
  mux2_1 U19959 ( .ip1(\LUT[97][12] ), .ip2(d[12]), .s(n17469), .op(n15030) );
  mux2_1 U19960 ( .ip1(\LUT[97][11] ), .ip2(d[11]), .s(n17469), .op(n15029) );
  mux2_1 U19961 ( .ip1(\LUT[97][10] ), .ip2(d[10]), .s(n17469), .op(n15028) );
  mux2_1 U19962 ( .ip1(\LUT[97][9] ), .ip2(d[9]), .s(n17469), .op(n15027) );
  mux2_1 U19963 ( .ip1(\LUT[97][8] ), .ip2(d[8]), .s(n17469), .op(n15026) );
  mux2_1 U19964 ( .ip1(\LUT[97][7] ), .ip2(d[7]), .s(n17469), .op(n15025) );
  mux2_1 U19965 ( .ip1(\LUT[97][6] ), .ip2(d[6]), .s(n17469), .op(n15024) );
  mux2_1 U19966 ( .ip1(\LUT[97][5] ), .ip2(d[5]), .s(n17470), .op(n15023) );
  mux2_1 U19967 ( .ip1(\LUT[97][4] ), .ip2(d[4]), .s(n17470), .op(n15022) );
  mux2_1 U19968 ( .ip1(\LUT[97][3] ), .ip2(d[3]), .s(n17470), .op(n15021) );
  mux2_1 U19969 ( .ip1(\LUT[97][2] ), .ip2(d[2]), .s(n17470), .op(n15020) );
  mux2_1 U19970 ( .ip1(\LUT[97][1] ), .ip2(d[1]), .s(n17470), .op(n15019) );
  mux2_1 U19971 ( .ip1(\LUT[97][0] ), .ip2(d[0]), .s(n17470), .op(n15018) );
  buf_1 U19972 ( .ip(d[15]), .op(n17541) );
  mux2_1 U19973 ( .ip1(\LUT[96][15] ), .ip2(n17541), .s(n17471), .op(n15017)
         );
  buf_1 U19974 ( .ip(d[14]), .op(n17542) );
  mux2_1 U19975 ( .ip1(\LUT[96][14] ), .ip2(n17542), .s(n17471), .op(n15016)
         );
  buf_1 U19976 ( .ip(d[13]), .op(n17543) );
  mux2_1 U19977 ( .ip1(\LUT[96][13] ), .ip2(n17543), .s(n17471), .op(n15015)
         );
  buf_1 U19978 ( .ip(d[12]), .op(n17544) );
  mux2_1 U19979 ( .ip1(\LUT[96][12] ), .ip2(n17544), .s(n17471), .op(n15014)
         );
  buf_1 U19980 ( .ip(d[11]), .op(n17545) );
  mux2_1 U19981 ( .ip1(\LUT[96][11] ), .ip2(n17545), .s(n17471), .op(n15013)
         );
  buf_1 U19982 ( .ip(d[10]), .op(n17546) );
  mux2_1 U19983 ( .ip1(\LUT[96][10] ), .ip2(n17546), .s(n17471), .op(n15012)
         );
  buf_1 U19984 ( .ip(d[9]), .op(n17547) );
  mux2_1 U19985 ( .ip1(\LUT[96][9] ), .ip2(n17547), .s(n17471), .op(n15011) );
  buf_1 U19986 ( .ip(d[8]), .op(n17548) );
  mux2_1 U19987 ( .ip1(\LUT[96][8] ), .ip2(n17548), .s(n17471), .op(n15010) );
  buf_1 U19988 ( .ip(d[7]), .op(n17549) );
  mux2_1 U19989 ( .ip1(\LUT[96][7] ), .ip2(n17549), .s(n17471), .op(n15009) );
  buf_1 U19990 ( .ip(d[6]), .op(n17551) );
  mux2_1 U19991 ( .ip1(\LUT[96][6] ), .ip2(n17551), .s(n17471), .op(n15008) );
  buf_1 U19992 ( .ip(d[5]), .op(n17552) );
  mux2_1 U19993 ( .ip1(\LUT[96][5] ), .ip2(n17552), .s(n17472), .op(n15007) );
  buf_1 U19994 ( .ip(d[4]), .op(n17553) );
  mux2_1 U19995 ( .ip1(\LUT[96][4] ), .ip2(n17553), .s(n17472), .op(n15006) );
  buf_1 U19996 ( .ip(d[3]), .op(n17554) );
  mux2_1 U19997 ( .ip1(\LUT[96][3] ), .ip2(n17554), .s(n17472), .op(n15005) );
  buf_1 U19998 ( .ip(d[2]), .op(n17555) );
  mux2_1 U19999 ( .ip1(\LUT[96][2] ), .ip2(n17555), .s(n17472), .op(n15004) );
  buf_1 U20000 ( .ip(d[1]), .op(n17556) );
  mux2_1 U20001 ( .ip1(\LUT[96][1] ), .ip2(n17556), .s(n17472), .op(n15003) );
  buf_1 U20002 ( .ip(d[0]), .op(n17558) );
  mux2_1 U20003 ( .ip1(\LUT[96][0] ), .ip2(n17558), .s(n17472), .op(n15002) );
  mux2_1 U20004 ( .ip1(\LUT[95][15] ), .ip2(n17541), .s(n17473), .op(n15001)
         );
  mux2_1 U20005 ( .ip1(\LUT[95][14] ), .ip2(n17542), .s(n17473), .op(n15000)
         );
  mux2_1 U20006 ( .ip1(\LUT[95][13] ), .ip2(n17543), .s(n17473), .op(n14999)
         );
  mux2_1 U20007 ( .ip1(\LUT[95][12] ), .ip2(n17544), .s(n17473), .op(n14998)
         );
  mux2_1 U20008 ( .ip1(\LUT[95][11] ), .ip2(n17545), .s(n17473), .op(n14997)
         );
  mux2_1 U20009 ( .ip1(\LUT[95][10] ), .ip2(n17546), .s(n17473), .op(n14996)
         );
  mux2_1 U20010 ( .ip1(\LUT[95][9] ), .ip2(n17547), .s(n17473), .op(n14995) );
  mux2_1 U20011 ( .ip1(\LUT[95][8] ), .ip2(n17548), .s(n17473), .op(n14994) );
  mux2_1 U20012 ( .ip1(\LUT[95][7] ), .ip2(n17549), .s(n17473), .op(n14993) );
  mux2_1 U20013 ( .ip1(\LUT[95][6] ), .ip2(n17551), .s(n17473), .op(n14992) );
  mux2_1 U20014 ( .ip1(\LUT[95][5] ), .ip2(n17552), .s(n17474), .op(n14991) );
  mux2_1 U20015 ( .ip1(\LUT[95][4] ), .ip2(n17553), .s(n17474), .op(n14990) );
  mux2_1 U20016 ( .ip1(\LUT[95][3] ), .ip2(n17554), .s(n17474), .op(n14989) );
  mux2_1 U20017 ( .ip1(\LUT[95][2] ), .ip2(n17555), .s(n17474), .op(n14988) );
  mux2_1 U20018 ( .ip1(\LUT[95][1] ), .ip2(n17556), .s(n17474), .op(n14987) );
  mux2_1 U20019 ( .ip1(\LUT[95][0] ), .ip2(n17558), .s(n17474), .op(n14986) );
  mux2_1 U20020 ( .ip1(\LUT[94][15] ), .ip2(n17541), .s(n17475), .op(n14985)
         );
  mux2_1 U20021 ( .ip1(\LUT[94][14] ), .ip2(n17542), .s(n17475), .op(n14984)
         );
  mux2_1 U20022 ( .ip1(\LUT[94][13] ), .ip2(n17543), .s(n17475), .op(n14983)
         );
  mux2_1 U20023 ( .ip1(\LUT[94][12] ), .ip2(n17544), .s(n17475), .op(n14982)
         );
  mux2_1 U20024 ( .ip1(\LUT[94][11] ), .ip2(n17545), .s(n17475), .op(n14981)
         );
  mux2_1 U20025 ( .ip1(\LUT[94][10] ), .ip2(n17546), .s(n17475), .op(n14980)
         );
  mux2_1 U20026 ( .ip1(\LUT[94][9] ), .ip2(n17547), .s(n17475), .op(n14979) );
  mux2_1 U20027 ( .ip1(\LUT[94][8] ), .ip2(n17548), .s(n17475), .op(n14978) );
  mux2_1 U20028 ( .ip1(\LUT[94][7] ), .ip2(n17549), .s(n17475), .op(n14977) );
  mux2_1 U20029 ( .ip1(\LUT[94][6] ), .ip2(n17551), .s(n17475), .op(n14976) );
  mux2_1 U20030 ( .ip1(\LUT[94][5] ), .ip2(n17552), .s(n17476), .op(n14975) );
  mux2_1 U20031 ( .ip1(\LUT[94][4] ), .ip2(n17553), .s(n17476), .op(n14974) );
  mux2_1 U20032 ( .ip1(\LUT[94][3] ), .ip2(n17554), .s(n17476), .op(n14973) );
  mux2_1 U20033 ( .ip1(\LUT[94][2] ), .ip2(n17555), .s(n17476), .op(n14972) );
  mux2_1 U20034 ( .ip1(\LUT[94][1] ), .ip2(n17556), .s(n17476), .op(n14971) );
  mux2_1 U20035 ( .ip1(\LUT[94][0] ), .ip2(n17558), .s(n17476), .op(n14970) );
  mux2_1 U20036 ( .ip1(\LUT[93][15] ), .ip2(n17541), .s(n17477), .op(n14969)
         );
  mux2_1 U20037 ( .ip1(\LUT[93][14] ), .ip2(n17542), .s(n17477), .op(n14968)
         );
  mux2_1 U20038 ( .ip1(\LUT[93][13] ), .ip2(n17543), .s(n17477), .op(n14967)
         );
  mux2_1 U20039 ( .ip1(\LUT[93][12] ), .ip2(n17544), .s(n17477), .op(n14966)
         );
  mux2_1 U20040 ( .ip1(\LUT[93][11] ), .ip2(n17545), .s(n17477), .op(n14965)
         );
  mux2_1 U20041 ( .ip1(\LUT[93][10] ), .ip2(n17546), .s(n17477), .op(n14964)
         );
  mux2_1 U20042 ( .ip1(\LUT[93][9] ), .ip2(n17547), .s(n17477), .op(n14963) );
  mux2_1 U20043 ( .ip1(\LUT[93][8] ), .ip2(n17548), .s(n17477), .op(n14962) );
  mux2_1 U20044 ( .ip1(\LUT[93][7] ), .ip2(n17549), .s(n17477), .op(n14961) );
  mux2_1 U20045 ( .ip1(\LUT[93][6] ), .ip2(n17551), .s(n17477), .op(n14960) );
  mux2_1 U20046 ( .ip1(\LUT[93][5] ), .ip2(n17552), .s(n17478), .op(n14959) );
  mux2_1 U20047 ( .ip1(\LUT[93][4] ), .ip2(n17553), .s(n17478), .op(n14958) );
  mux2_1 U20048 ( .ip1(\LUT[93][3] ), .ip2(n17554), .s(n17478), .op(n14957) );
  mux2_1 U20049 ( .ip1(\LUT[93][2] ), .ip2(n17555), .s(n17478), .op(n14956) );
  mux2_1 U20050 ( .ip1(\LUT[93][1] ), .ip2(n17556), .s(n17478), .op(n14955) );
  mux2_1 U20051 ( .ip1(\LUT[93][0] ), .ip2(n17558), .s(n17478), .op(n14954) );
  mux2_1 U20052 ( .ip1(\LUT[92][15] ), .ip2(n17541), .s(n17479), .op(n14953)
         );
  mux2_1 U20053 ( .ip1(\LUT[92][14] ), .ip2(n17542), .s(n17479), .op(n14952)
         );
  mux2_1 U20054 ( .ip1(\LUT[92][13] ), .ip2(n17543), .s(n17479), .op(n14951)
         );
  mux2_1 U20055 ( .ip1(\LUT[92][12] ), .ip2(n17544), .s(n17479), .op(n14950)
         );
  mux2_1 U20056 ( .ip1(\LUT[92][11] ), .ip2(n17545), .s(n17479), .op(n14949)
         );
  mux2_1 U20057 ( .ip1(\LUT[92][10] ), .ip2(n17546), .s(n17479), .op(n14948)
         );
  mux2_1 U20058 ( .ip1(\LUT[92][9] ), .ip2(n17547), .s(n17479), .op(n14947) );
  mux2_1 U20059 ( .ip1(\LUT[92][8] ), .ip2(n17548), .s(n17479), .op(n14946) );
  mux2_1 U20060 ( .ip1(\LUT[92][7] ), .ip2(n17549), .s(n17479), .op(n14945) );
  mux2_1 U20061 ( .ip1(\LUT[92][6] ), .ip2(n17551), .s(n17479), .op(n14944) );
  mux2_1 U20062 ( .ip1(\LUT[92][5] ), .ip2(n17552), .s(n17480), .op(n14943) );
  mux2_1 U20063 ( .ip1(\LUT[92][4] ), .ip2(n17553), .s(n17480), .op(n14942) );
  mux2_1 U20064 ( .ip1(\LUT[92][3] ), .ip2(n17554), .s(n17480), .op(n14941) );
  mux2_1 U20065 ( .ip1(\LUT[92][2] ), .ip2(n17555), .s(n17480), .op(n14940) );
  mux2_1 U20066 ( .ip1(\LUT[92][1] ), .ip2(n17556), .s(n17480), .op(n14939) );
  mux2_1 U20067 ( .ip1(\LUT[92][0] ), .ip2(n17558), .s(n17480), .op(n14938) );
  mux2_1 U20068 ( .ip1(\LUT[91][15] ), .ip2(n17541), .s(n17481), .op(n14937)
         );
  mux2_1 U20069 ( .ip1(\LUT[91][14] ), .ip2(n17542), .s(n17481), .op(n14936)
         );
  mux2_1 U20070 ( .ip1(\LUT[91][13] ), .ip2(n17543), .s(n17481), .op(n14935)
         );
  mux2_1 U20071 ( .ip1(\LUT[91][12] ), .ip2(n17544), .s(n17481), .op(n14934)
         );
  mux2_1 U20072 ( .ip1(\LUT[91][11] ), .ip2(n17545), .s(n17481), .op(n14933)
         );
  mux2_1 U20073 ( .ip1(\LUT[91][10] ), .ip2(n17546), .s(n17481), .op(n14932)
         );
  mux2_1 U20074 ( .ip1(\LUT[91][9] ), .ip2(n17547), .s(n17481), .op(n14931) );
  mux2_1 U20075 ( .ip1(\LUT[91][8] ), .ip2(n17548), .s(n17481), .op(n14930) );
  mux2_1 U20076 ( .ip1(\LUT[91][7] ), .ip2(n17549), .s(n17481), .op(n14929) );
  mux2_1 U20077 ( .ip1(\LUT[91][6] ), .ip2(n17551), .s(n17481), .op(n14928) );
  mux2_1 U20078 ( .ip1(\LUT[91][5] ), .ip2(n17552), .s(n17482), .op(n14927) );
  mux2_1 U20079 ( .ip1(\LUT[91][4] ), .ip2(n17553), .s(n17482), .op(n14926) );
  mux2_1 U20080 ( .ip1(\LUT[91][3] ), .ip2(n17554), .s(n17482), .op(n14925) );
  mux2_1 U20081 ( .ip1(\LUT[91][2] ), .ip2(n17555), .s(n17482), .op(n14924) );
  mux2_1 U20082 ( .ip1(\LUT[91][1] ), .ip2(n17556), .s(n17482), .op(n14923) );
  mux2_1 U20083 ( .ip1(\LUT[91][0] ), .ip2(n17558), .s(n17482), .op(n14922) );
  mux2_1 U20084 ( .ip1(\LUT[90][15] ), .ip2(n17541), .s(n17483), .op(n14921)
         );
  mux2_1 U20085 ( .ip1(\LUT[90][14] ), .ip2(n17542), .s(n17483), .op(n14920)
         );
  mux2_1 U20086 ( .ip1(\LUT[90][13] ), .ip2(n17543), .s(n17483), .op(n14919)
         );
  mux2_1 U20087 ( .ip1(\LUT[90][12] ), .ip2(n17544), .s(n17483), .op(n14918)
         );
  mux2_1 U20088 ( .ip1(\LUT[90][11] ), .ip2(n17545), .s(n17483), .op(n14917)
         );
  mux2_1 U20089 ( .ip1(\LUT[90][10] ), .ip2(n17546), .s(n17483), .op(n14916)
         );
  mux2_1 U20090 ( .ip1(\LUT[90][9] ), .ip2(n17547), .s(n17483), .op(n14915) );
  mux2_1 U20091 ( .ip1(\LUT[90][8] ), .ip2(n17548), .s(n17483), .op(n14914) );
  mux2_1 U20092 ( .ip1(\LUT[90][7] ), .ip2(n17549), .s(n17483), .op(n14913) );
  mux2_1 U20093 ( .ip1(\LUT[90][6] ), .ip2(n17551), .s(n17483), .op(n14912) );
  mux2_1 U20094 ( .ip1(\LUT[90][5] ), .ip2(n17552), .s(n17484), .op(n14911) );
  mux2_1 U20095 ( .ip1(\LUT[90][4] ), .ip2(n17553), .s(n17484), .op(n14910) );
  mux2_1 U20096 ( .ip1(\LUT[90][3] ), .ip2(n17554), .s(n17484), .op(n14909) );
  mux2_1 U20097 ( .ip1(\LUT[90][2] ), .ip2(n17555), .s(n17484), .op(n14908) );
  mux2_1 U20098 ( .ip1(\LUT[90][1] ), .ip2(n17556), .s(n17484), .op(n14907) );
  mux2_1 U20099 ( .ip1(\LUT[90][0] ), .ip2(n17558), .s(n17484), .op(n14906) );
  mux2_1 U20100 ( .ip1(\LUT[89][15] ), .ip2(n17541), .s(n17485), .op(n14905)
         );
  mux2_1 U20101 ( .ip1(\LUT[89][14] ), .ip2(n17542), .s(n17485), .op(n14904)
         );
  mux2_1 U20102 ( .ip1(\LUT[89][13] ), .ip2(n17543), .s(n17485), .op(n14903)
         );
  mux2_1 U20103 ( .ip1(\LUT[89][12] ), .ip2(n17544), .s(n17485), .op(n14902)
         );
  mux2_1 U20104 ( .ip1(\LUT[89][11] ), .ip2(n17545), .s(n17485), .op(n14901)
         );
  mux2_1 U20105 ( .ip1(\LUT[89][10] ), .ip2(n17546), .s(n17485), .op(n14900)
         );
  mux2_1 U20106 ( .ip1(\LUT[89][9] ), .ip2(n17547), .s(n17485), .op(n14899) );
  mux2_1 U20107 ( .ip1(\LUT[89][8] ), .ip2(n17548), .s(n17485), .op(n14898) );
  mux2_1 U20108 ( .ip1(\LUT[89][7] ), .ip2(n17549), .s(n17485), .op(n14897) );
  mux2_1 U20109 ( .ip1(\LUT[89][6] ), .ip2(n17551), .s(n17485), .op(n14896) );
  mux2_1 U20110 ( .ip1(\LUT[89][5] ), .ip2(n17552), .s(n17486), .op(n14895) );
  mux2_1 U20111 ( .ip1(\LUT[89][4] ), .ip2(n17553), .s(n17486), .op(n14894) );
  mux2_1 U20112 ( .ip1(\LUT[89][3] ), .ip2(n17554), .s(n17486), .op(n14893) );
  mux2_1 U20113 ( .ip1(\LUT[89][2] ), .ip2(n17555), .s(n17486), .op(n14892) );
  mux2_1 U20114 ( .ip1(\LUT[89][1] ), .ip2(n17556), .s(n17486), .op(n14891) );
  mux2_1 U20115 ( .ip1(\LUT[89][0] ), .ip2(n17558), .s(n17486), .op(n14890) );
  mux2_1 U20116 ( .ip1(\LUT[88][15] ), .ip2(n17541), .s(n17487), .op(n14889)
         );
  mux2_1 U20117 ( .ip1(\LUT[88][14] ), .ip2(n17542), .s(n17487), .op(n14888)
         );
  mux2_1 U20118 ( .ip1(\LUT[88][13] ), .ip2(n17543), .s(n17487), .op(n14887)
         );
  mux2_1 U20119 ( .ip1(\LUT[88][12] ), .ip2(n17544), .s(n17487), .op(n14886)
         );
  mux2_1 U20120 ( .ip1(\LUT[88][11] ), .ip2(n17545), .s(n17487), .op(n14885)
         );
  mux2_1 U20121 ( .ip1(\LUT[88][10] ), .ip2(n17546), .s(n17487), .op(n14884)
         );
  mux2_1 U20122 ( .ip1(\LUT[88][9] ), .ip2(n17547), .s(n17487), .op(n14883) );
  mux2_1 U20123 ( .ip1(\LUT[88][8] ), .ip2(n17548), .s(n17487), .op(n14882) );
  mux2_1 U20124 ( .ip1(\LUT[88][7] ), .ip2(n17549), .s(n17487), .op(n14881) );
  mux2_1 U20125 ( .ip1(\LUT[88][6] ), .ip2(n17551), .s(n17487), .op(n14880) );
  mux2_1 U20126 ( .ip1(\LUT[88][5] ), .ip2(n17552), .s(n17488), .op(n14879) );
  mux2_1 U20127 ( .ip1(\LUT[88][4] ), .ip2(n17553), .s(n17488), .op(n14878) );
  mux2_1 U20128 ( .ip1(\LUT[88][3] ), .ip2(n17554), .s(n17488), .op(n14877) );
  mux2_1 U20129 ( .ip1(\LUT[88][2] ), .ip2(n17555), .s(n17488), .op(n14876) );
  mux2_1 U20130 ( .ip1(\LUT[88][1] ), .ip2(n17556), .s(n17488), .op(n14875) );
  mux2_1 U20131 ( .ip1(\LUT[88][0] ), .ip2(n17558), .s(n17488), .op(n14874) );
  mux2_1 U20132 ( .ip1(\LUT[87][15] ), .ip2(n17541), .s(n17489), .op(n14873)
         );
  mux2_1 U20133 ( .ip1(\LUT[87][14] ), .ip2(n17542), .s(n17489), .op(n14872)
         );
  mux2_1 U20134 ( .ip1(\LUT[87][13] ), .ip2(n17543), .s(n17489), .op(n14871)
         );
  mux2_1 U20135 ( .ip1(\LUT[87][12] ), .ip2(n17544), .s(n17489), .op(n14870)
         );
  mux2_1 U20136 ( .ip1(\LUT[87][11] ), .ip2(n17545), .s(n17489), .op(n14869)
         );
  mux2_1 U20137 ( .ip1(\LUT[87][10] ), .ip2(n17546), .s(n17489), .op(n14868)
         );
  mux2_1 U20138 ( .ip1(\LUT[87][9] ), .ip2(n17547), .s(n17489), .op(n14867) );
  mux2_1 U20139 ( .ip1(\LUT[87][8] ), .ip2(n17548), .s(n17489), .op(n14866) );
  mux2_1 U20140 ( .ip1(\LUT[87][7] ), .ip2(n17549), .s(n17489), .op(n14865) );
  mux2_1 U20141 ( .ip1(\LUT[87][6] ), .ip2(n17551), .s(n17489), .op(n14864) );
  mux2_1 U20142 ( .ip1(\LUT[87][5] ), .ip2(n17552), .s(n17490), .op(n14863) );
  mux2_1 U20143 ( .ip1(\LUT[87][4] ), .ip2(n17553), .s(n17490), .op(n14862) );
  mux2_1 U20144 ( .ip1(\LUT[87][3] ), .ip2(n17554), .s(n17490), .op(n14861) );
  mux2_1 U20145 ( .ip1(\LUT[87][2] ), .ip2(n17555), .s(n17490), .op(n14860) );
  mux2_1 U20146 ( .ip1(\LUT[87][1] ), .ip2(n17556), .s(n17490), .op(n14859) );
  mux2_1 U20147 ( .ip1(\LUT[87][0] ), .ip2(n17558), .s(n17490), .op(n14858) );
  mux2_1 U20148 ( .ip1(\LUT[86][15] ), .ip2(n17541), .s(n17491), .op(n14857)
         );
  mux2_1 U20149 ( .ip1(\LUT[86][14] ), .ip2(n17542), .s(n17491), .op(n14856)
         );
  mux2_1 U20150 ( .ip1(\LUT[86][13] ), .ip2(n17543), .s(n17491), .op(n14855)
         );
  mux2_1 U20151 ( .ip1(\LUT[86][12] ), .ip2(n17544), .s(n17491), .op(n14854)
         );
  mux2_1 U20152 ( .ip1(\LUT[86][11] ), .ip2(n17545), .s(n17491), .op(n14853)
         );
  mux2_1 U20153 ( .ip1(\LUT[86][10] ), .ip2(n17546), .s(n17491), .op(n14852)
         );
  mux2_1 U20154 ( .ip1(\LUT[86][9] ), .ip2(n17547), .s(n17491), .op(n14851) );
  mux2_1 U20155 ( .ip1(\LUT[86][8] ), .ip2(n17548), .s(n17491), .op(n14850) );
  mux2_1 U20156 ( .ip1(\LUT[86][7] ), .ip2(n17549), .s(n17491), .op(n14849) );
  mux2_1 U20157 ( .ip1(\LUT[86][6] ), .ip2(n17551), .s(n17491), .op(n14848) );
  mux2_1 U20158 ( .ip1(\LUT[86][5] ), .ip2(n17552), .s(n17492), .op(n14847) );
  mux2_1 U20159 ( .ip1(\LUT[86][4] ), .ip2(n17553), .s(n17492), .op(n14846) );
  mux2_1 U20160 ( .ip1(\LUT[86][3] ), .ip2(n17554), .s(n17492), .op(n14845) );
  mux2_1 U20161 ( .ip1(\LUT[86][2] ), .ip2(n17555), .s(n17492), .op(n14844) );
  mux2_1 U20162 ( .ip1(\LUT[86][1] ), .ip2(n17556), .s(n17492), .op(n14843) );
  mux2_1 U20163 ( .ip1(\LUT[86][0] ), .ip2(n17558), .s(n17492), .op(n14842) );
  mux2_1 U20164 ( .ip1(\LUT[85][15] ), .ip2(n17541), .s(n17493), .op(n14841)
         );
  mux2_1 U20165 ( .ip1(\LUT[85][14] ), .ip2(n17542), .s(n17493), .op(n14840)
         );
  mux2_1 U20166 ( .ip1(\LUT[85][13] ), .ip2(n17543), .s(n17493), .op(n14839)
         );
  mux2_1 U20167 ( .ip1(\LUT[85][12] ), .ip2(n17544), .s(n17493), .op(n14838)
         );
  mux2_1 U20168 ( .ip1(\LUT[85][11] ), .ip2(n17545), .s(n17493), .op(n14837)
         );
  mux2_1 U20169 ( .ip1(\LUT[85][10] ), .ip2(n17546), .s(n17493), .op(n14836)
         );
  mux2_1 U20170 ( .ip1(\LUT[85][9] ), .ip2(n17547), .s(n17493), .op(n14835) );
  mux2_1 U20171 ( .ip1(\LUT[85][8] ), .ip2(n17548), .s(n17493), .op(n14834) );
  mux2_1 U20172 ( .ip1(\LUT[85][7] ), .ip2(n17549), .s(n17493), .op(n14833) );
  mux2_1 U20173 ( .ip1(\LUT[85][6] ), .ip2(n17551), .s(n17493), .op(n14832) );
  mux2_1 U20174 ( .ip1(\LUT[85][5] ), .ip2(n17552), .s(n17494), .op(n14831) );
  mux2_1 U20175 ( .ip1(\LUT[85][4] ), .ip2(n17553), .s(n17494), .op(n14830) );
  mux2_1 U20176 ( .ip1(\LUT[85][3] ), .ip2(n17554), .s(n17494), .op(n14829) );
  mux2_1 U20177 ( .ip1(\LUT[85][2] ), .ip2(n17555), .s(n17494), .op(n14828) );
  mux2_1 U20178 ( .ip1(\LUT[85][1] ), .ip2(n17556), .s(n17494), .op(n14827) );
  mux2_1 U20179 ( .ip1(\LUT[85][0] ), .ip2(n17558), .s(n17494), .op(n14826) );
  mux2_1 U20180 ( .ip1(\LUT[84][15] ), .ip2(n17541), .s(n17495), .op(n14825)
         );
  mux2_1 U20181 ( .ip1(\LUT[84][14] ), .ip2(n17542), .s(n17495), .op(n14824)
         );
  mux2_1 U20182 ( .ip1(\LUT[84][13] ), .ip2(n17543), .s(n17495), .op(n14823)
         );
  mux2_1 U20183 ( .ip1(\LUT[84][12] ), .ip2(n17544), .s(n17495), .op(n14822)
         );
  mux2_1 U20184 ( .ip1(\LUT[84][11] ), .ip2(n17545), .s(n17495), .op(n14821)
         );
  mux2_1 U20185 ( .ip1(\LUT[84][10] ), .ip2(n17546), .s(n17495), .op(n14820)
         );
  mux2_1 U20186 ( .ip1(\LUT[84][9] ), .ip2(n17547), .s(n17495), .op(n14819) );
  mux2_1 U20187 ( .ip1(\LUT[84][8] ), .ip2(n17548), .s(n17495), .op(n14818) );
  mux2_1 U20188 ( .ip1(\LUT[84][7] ), .ip2(n17549), .s(n17495), .op(n14817) );
  mux2_1 U20189 ( .ip1(\LUT[84][6] ), .ip2(n17551), .s(n17495), .op(n14816) );
  mux2_1 U20190 ( .ip1(\LUT[84][5] ), .ip2(n17552), .s(n17496), .op(n14815) );
  mux2_1 U20191 ( .ip1(\LUT[84][4] ), .ip2(n17553), .s(n17496), .op(n14814) );
  mux2_1 U20192 ( .ip1(\LUT[84][3] ), .ip2(n17554), .s(n17496), .op(n14813) );
  mux2_1 U20193 ( .ip1(\LUT[84][2] ), .ip2(n17555), .s(n17496), .op(n14812) );
  mux2_1 U20194 ( .ip1(\LUT[84][1] ), .ip2(n17556), .s(n17496), .op(n14811) );
  mux2_1 U20195 ( .ip1(\LUT[84][0] ), .ip2(n17558), .s(n17496), .op(n14810) );
  mux2_1 U20196 ( .ip1(\LUT[83][15] ), .ip2(n17541), .s(n17497), .op(n14809)
         );
  mux2_1 U20197 ( .ip1(\LUT[83][14] ), .ip2(n17542), .s(n17497), .op(n14808)
         );
  mux2_1 U20198 ( .ip1(\LUT[83][13] ), .ip2(n17543), .s(n17497), .op(n14807)
         );
  mux2_1 U20199 ( .ip1(\LUT[83][12] ), .ip2(n17544), .s(n17497), .op(n14806)
         );
  mux2_1 U20200 ( .ip1(\LUT[83][11] ), .ip2(n17545), .s(n17497), .op(n14805)
         );
  mux2_1 U20201 ( .ip1(\LUT[83][10] ), .ip2(n17546), .s(n17497), .op(n14804)
         );
  mux2_1 U20202 ( .ip1(\LUT[83][9] ), .ip2(n17547), .s(n17497), .op(n14803) );
  mux2_1 U20203 ( .ip1(\LUT[83][8] ), .ip2(n17548), .s(n17497), .op(n14802) );
  mux2_1 U20204 ( .ip1(\LUT[83][7] ), .ip2(n17549), .s(n17497), .op(n14801) );
  mux2_1 U20205 ( .ip1(\LUT[83][6] ), .ip2(n17551), .s(n17497), .op(n14800) );
  mux2_1 U20206 ( .ip1(\LUT[83][5] ), .ip2(n17552), .s(n17498), .op(n14799) );
  mux2_1 U20207 ( .ip1(\LUT[83][4] ), .ip2(n17553), .s(n17498), .op(n14798) );
  mux2_1 U20208 ( .ip1(\LUT[83][3] ), .ip2(n17554), .s(n17498), .op(n14797) );
  mux2_1 U20209 ( .ip1(\LUT[83][2] ), .ip2(n17555), .s(n17498), .op(n14796) );
  mux2_1 U20210 ( .ip1(\LUT[83][1] ), .ip2(n17556), .s(n17498), .op(n14795) );
  mux2_1 U20211 ( .ip1(\LUT[83][0] ), .ip2(n17558), .s(n17498), .op(n14794) );
  mux2_1 U20212 ( .ip1(\LUT[82][15] ), .ip2(n17541), .s(n17499), .op(n14793)
         );
  mux2_1 U20213 ( .ip1(\LUT[82][14] ), .ip2(n17542), .s(n17499), .op(n14792)
         );
  mux2_1 U20214 ( .ip1(\LUT[82][13] ), .ip2(n17543), .s(n17499), .op(n14791)
         );
  mux2_1 U20215 ( .ip1(\LUT[82][12] ), .ip2(n17544), .s(n17499), .op(n14790)
         );
  mux2_1 U20216 ( .ip1(\LUT[82][11] ), .ip2(n17545), .s(n17499), .op(n14789)
         );
  mux2_1 U20217 ( .ip1(\LUT[82][10] ), .ip2(n17546), .s(n17499), .op(n14788)
         );
  mux2_1 U20218 ( .ip1(\LUT[82][9] ), .ip2(n17547), .s(n17499), .op(n14787) );
  mux2_1 U20219 ( .ip1(\LUT[82][8] ), .ip2(n17548), .s(n17499), .op(n14786) );
  mux2_1 U20220 ( .ip1(\LUT[82][7] ), .ip2(n17549), .s(n17499), .op(n14785) );
  mux2_1 U20221 ( .ip1(\LUT[82][6] ), .ip2(n17551), .s(n17499), .op(n14784) );
  mux2_1 U20222 ( .ip1(\LUT[82][5] ), .ip2(n17552), .s(n17500), .op(n14783) );
  mux2_1 U20223 ( .ip1(\LUT[82][4] ), .ip2(n17553), .s(n17500), .op(n14782) );
  mux2_1 U20224 ( .ip1(\LUT[82][3] ), .ip2(n17554), .s(n17500), .op(n14781) );
  mux2_1 U20225 ( .ip1(\LUT[82][2] ), .ip2(n17555), .s(n17500), .op(n14780) );
  mux2_1 U20226 ( .ip1(\LUT[82][1] ), .ip2(n17556), .s(n17500), .op(n14779) );
  mux2_1 U20227 ( .ip1(\LUT[82][0] ), .ip2(n17558), .s(n17500), .op(n14778) );
  mux2_1 U20228 ( .ip1(\LUT[81][15] ), .ip2(n17541), .s(n17501), .op(n14777)
         );
  mux2_1 U20229 ( .ip1(\LUT[81][14] ), .ip2(n17542), .s(n17501), .op(n14776)
         );
  mux2_1 U20230 ( .ip1(\LUT[81][13] ), .ip2(n17543), .s(n17501), .op(n14775)
         );
  mux2_1 U20231 ( .ip1(\LUT[81][12] ), .ip2(n17544), .s(n17501), .op(n14774)
         );
  mux2_1 U20232 ( .ip1(\LUT[81][11] ), .ip2(n17545), .s(n17501), .op(n14773)
         );
  mux2_1 U20233 ( .ip1(\LUT[81][10] ), .ip2(n17546), .s(n17501), .op(n14772)
         );
  mux2_1 U20234 ( .ip1(\LUT[81][9] ), .ip2(n17547), .s(n17501), .op(n14771) );
  mux2_1 U20235 ( .ip1(\LUT[81][8] ), .ip2(n17548), .s(n17501), .op(n14770) );
  mux2_1 U20236 ( .ip1(\LUT[81][7] ), .ip2(n17549), .s(n17501), .op(n14769) );
  mux2_1 U20237 ( .ip1(\LUT[81][6] ), .ip2(n17551), .s(n17501), .op(n14768) );
  mux2_1 U20238 ( .ip1(\LUT[81][5] ), .ip2(n17552), .s(n17502), .op(n14767) );
  mux2_1 U20239 ( .ip1(\LUT[81][4] ), .ip2(n17553), .s(n17502), .op(n14766) );
  mux2_1 U20240 ( .ip1(\LUT[81][3] ), .ip2(n17554), .s(n17502), .op(n14765) );
  mux2_1 U20241 ( .ip1(\LUT[81][2] ), .ip2(n17555), .s(n17502), .op(n14764) );
  mux2_1 U20242 ( .ip1(\LUT[81][1] ), .ip2(n17556), .s(n17502), .op(n14763) );
  mux2_1 U20243 ( .ip1(\LUT[81][0] ), .ip2(n17558), .s(n17502), .op(n14762) );
  mux2_1 U20244 ( .ip1(\LUT[80][15] ), .ip2(n17541), .s(n17503), .op(n14761)
         );
  mux2_1 U20245 ( .ip1(\LUT[80][14] ), .ip2(n17542), .s(n17503), .op(n14760)
         );
  mux2_1 U20246 ( .ip1(\LUT[80][13] ), .ip2(n17543), .s(n17503), .op(n14759)
         );
  mux2_1 U20247 ( .ip1(\LUT[80][12] ), .ip2(n17544), .s(n17503), .op(n14758)
         );
  mux2_1 U20248 ( .ip1(\LUT[80][11] ), .ip2(n17545), .s(n17503), .op(n14757)
         );
  mux2_1 U20249 ( .ip1(\LUT[80][10] ), .ip2(n17546), .s(n17503), .op(n14756)
         );
  mux2_1 U20250 ( .ip1(\LUT[80][9] ), .ip2(n17547), .s(n17503), .op(n14755) );
  mux2_1 U20251 ( .ip1(\LUT[80][8] ), .ip2(n17548), .s(n17503), .op(n14754) );
  mux2_1 U20252 ( .ip1(\LUT[80][7] ), .ip2(n17549), .s(n17503), .op(n14753) );
  mux2_1 U20253 ( .ip1(\LUT[80][6] ), .ip2(n17551), .s(n17503), .op(n14752) );
  mux2_1 U20254 ( .ip1(\LUT[80][5] ), .ip2(n17552), .s(n17504), .op(n14751) );
  mux2_1 U20255 ( .ip1(\LUT[80][4] ), .ip2(n17553), .s(n17504), .op(n14750) );
  mux2_1 U20256 ( .ip1(\LUT[80][3] ), .ip2(n17554), .s(n17504), .op(n14749) );
  mux2_1 U20257 ( .ip1(\LUT[80][2] ), .ip2(n17555), .s(n17504), .op(n14748) );
  mux2_1 U20258 ( .ip1(\LUT[80][1] ), .ip2(n17556), .s(n17504), .op(n14747) );
  mux2_1 U20259 ( .ip1(\LUT[80][0] ), .ip2(n17558), .s(n17504), .op(n14746) );
  mux2_1 U20260 ( .ip1(\LUT[79][15] ), .ip2(n17541), .s(n17505), .op(n14745)
         );
  mux2_1 U20261 ( .ip1(\LUT[79][14] ), .ip2(n17542), .s(n17505), .op(n14744)
         );
  mux2_1 U20262 ( .ip1(\LUT[79][13] ), .ip2(n17543), .s(n17505), .op(n14743)
         );
  mux2_1 U20263 ( .ip1(\LUT[79][12] ), .ip2(n17544), .s(n17505), .op(n14742)
         );
  mux2_1 U20264 ( .ip1(\LUT[79][11] ), .ip2(n17545), .s(n17505), .op(n14741)
         );
  mux2_1 U20265 ( .ip1(\LUT[79][10] ), .ip2(n17546), .s(n17505), .op(n14740)
         );
  mux2_1 U20266 ( .ip1(\LUT[79][9] ), .ip2(n17547), .s(n17505), .op(n14739) );
  mux2_1 U20267 ( .ip1(\LUT[79][8] ), .ip2(n17548), .s(n17505), .op(n14738) );
  mux2_1 U20268 ( .ip1(\LUT[79][7] ), .ip2(n17549), .s(n17505), .op(n14737) );
  mux2_1 U20269 ( .ip1(\LUT[79][6] ), .ip2(n17551), .s(n17505), .op(n14736) );
  mux2_1 U20270 ( .ip1(\LUT[79][5] ), .ip2(n17552), .s(n17506), .op(n14735) );
  mux2_1 U20271 ( .ip1(\LUT[79][4] ), .ip2(n17553), .s(n17506), .op(n14734) );
  mux2_1 U20272 ( .ip1(\LUT[79][3] ), .ip2(n17554), .s(n17506), .op(n14733) );
  mux2_1 U20273 ( .ip1(\LUT[79][2] ), .ip2(n17555), .s(n17506), .op(n14732) );
  mux2_1 U20274 ( .ip1(\LUT[79][1] ), .ip2(n17556), .s(n17506), .op(n14731) );
  mux2_1 U20275 ( .ip1(\LUT[79][0] ), .ip2(n17558), .s(n17506), .op(n14730) );
  mux2_1 U20276 ( .ip1(\LUT[78][15] ), .ip2(n17541), .s(n17507), .op(n14729)
         );
  mux2_1 U20277 ( .ip1(\LUT[78][14] ), .ip2(n17542), .s(n17507), .op(n14728)
         );
  mux2_1 U20278 ( .ip1(\LUT[78][13] ), .ip2(n17543), .s(n17507), .op(n14727)
         );
  mux2_1 U20279 ( .ip1(\LUT[78][12] ), .ip2(n17544), .s(n17507), .op(n14726)
         );
  mux2_1 U20280 ( .ip1(\LUT[78][11] ), .ip2(n17545), .s(n17507), .op(n14725)
         );
  mux2_1 U20281 ( .ip1(\LUT[78][10] ), .ip2(n17546), .s(n17507), .op(n14724)
         );
  mux2_1 U20282 ( .ip1(\LUT[78][9] ), .ip2(n17547), .s(n17507), .op(n14723) );
  mux2_1 U20283 ( .ip1(\LUT[78][8] ), .ip2(n17548), .s(n17507), .op(n14722) );
  mux2_1 U20284 ( .ip1(\LUT[78][7] ), .ip2(n17549), .s(n17507), .op(n14721) );
  mux2_1 U20285 ( .ip1(\LUT[78][6] ), .ip2(n17551), .s(n17507), .op(n14720) );
  mux2_1 U20286 ( .ip1(\LUT[78][5] ), .ip2(n17552), .s(n17508), .op(n14719) );
  mux2_1 U20287 ( .ip1(\LUT[78][4] ), .ip2(n17553), .s(n17508), .op(n14718) );
  mux2_1 U20288 ( .ip1(\LUT[78][3] ), .ip2(n17554), .s(n17508), .op(n14717) );
  mux2_1 U20289 ( .ip1(\LUT[78][2] ), .ip2(n17555), .s(n17508), .op(n14716) );
  mux2_1 U20290 ( .ip1(\LUT[78][1] ), .ip2(n17556), .s(n17508), .op(n14715) );
  mux2_1 U20291 ( .ip1(\LUT[78][0] ), .ip2(n17558), .s(n17508), .op(n14714) );
  mux2_1 U20292 ( .ip1(\LUT[77][15] ), .ip2(n17541), .s(n17509), .op(n14713)
         );
  mux2_1 U20293 ( .ip1(\LUT[77][14] ), .ip2(n17542), .s(n17509), .op(n14712)
         );
  mux2_1 U20294 ( .ip1(\LUT[77][13] ), .ip2(n17543), .s(n17509), .op(n14711)
         );
  mux2_1 U20295 ( .ip1(\LUT[77][12] ), .ip2(n17544), .s(n17509), .op(n14710)
         );
  mux2_1 U20296 ( .ip1(\LUT[77][11] ), .ip2(n17545), .s(n17509), .op(n14709)
         );
  mux2_1 U20297 ( .ip1(\LUT[77][10] ), .ip2(n17546), .s(n17509), .op(n14708)
         );
  mux2_1 U20298 ( .ip1(\LUT[77][9] ), .ip2(n17547), .s(n17509), .op(n14707) );
  mux2_1 U20299 ( .ip1(\LUT[77][8] ), .ip2(n17548), .s(n17509), .op(n14706) );
  mux2_1 U20300 ( .ip1(\LUT[77][7] ), .ip2(n17549), .s(n17509), .op(n14705) );
  mux2_1 U20301 ( .ip1(\LUT[77][6] ), .ip2(n17551), .s(n17509), .op(n14704) );
  mux2_1 U20302 ( .ip1(\LUT[77][5] ), .ip2(n17552), .s(n17510), .op(n14703) );
  mux2_1 U20303 ( .ip1(\LUT[77][4] ), .ip2(n17553), .s(n17510), .op(n14702) );
  mux2_1 U20304 ( .ip1(\LUT[77][3] ), .ip2(n17554), .s(n17510), .op(n14701) );
  mux2_1 U20305 ( .ip1(\LUT[77][2] ), .ip2(n17555), .s(n17510), .op(n14700) );
  mux2_1 U20306 ( .ip1(\LUT[77][1] ), .ip2(n17556), .s(n17510), .op(n14699) );
  mux2_1 U20307 ( .ip1(\LUT[77][0] ), .ip2(n17558), .s(n17510), .op(n14698) );
  mux2_1 U20308 ( .ip1(\LUT[76][15] ), .ip2(n17541), .s(n17511), .op(n14697)
         );
  mux2_1 U20309 ( .ip1(\LUT[76][14] ), .ip2(n17542), .s(n17511), .op(n14696)
         );
  mux2_1 U20310 ( .ip1(\LUT[76][13] ), .ip2(n17543), .s(n17511), .op(n14695)
         );
  mux2_1 U20311 ( .ip1(\LUT[76][12] ), .ip2(n17544), .s(n17511), .op(n14694)
         );
  mux2_1 U20312 ( .ip1(\LUT[76][11] ), .ip2(n17545), .s(n17511), .op(n14693)
         );
  mux2_1 U20313 ( .ip1(\LUT[76][10] ), .ip2(n17546), .s(n17511), .op(n14692)
         );
  mux2_1 U20314 ( .ip1(\LUT[76][9] ), .ip2(n17547), .s(n17511), .op(n14691) );
  mux2_1 U20315 ( .ip1(\LUT[76][8] ), .ip2(n17548), .s(n17511), .op(n14690) );
  mux2_1 U20316 ( .ip1(\LUT[76][7] ), .ip2(n17549), .s(n17511), .op(n14689) );
  mux2_1 U20317 ( .ip1(\LUT[76][6] ), .ip2(n17551), .s(n17511), .op(n14688) );
  mux2_1 U20318 ( .ip1(\LUT[76][5] ), .ip2(n17552), .s(n17512), .op(n14687) );
  mux2_1 U20319 ( .ip1(\LUT[76][4] ), .ip2(n17553), .s(n17512), .op(n14686) );
  mux2_1 U20320 ( .ip1(\LUT[76][3] ), .ip2(n17554), .s(n17512), .op(n14685) );
  mux2_1 U20321 ( .ip1(\LUT[76][2] ), .ip2(n17555), .s(n17512), .op(n14684) );
  mux2_1 U20322 ( .ip1(\LUT[76][1] ), .ip2(n17556), .s(n17512), .op(n14683) );
  mux2_1 U20323 ( .ip1(\LUT[76][0] ), .ip2(n17558), .s(n17512), .op(n14682) );
  mux2_1 U20324 ( .ip1(\LUT[75][15] ), .ip2(n17541), .s(n17513), .op(n14681)
         );
  mux2_1 U20325 ( .ip1(\LUT[75][14] ), .ip2(n17542), .s(n17513), .op(n14680)
         );
  mux2_1 U20326 ( .ip1(\LUT[75][13] ), .ip2(n17543), .s(n17513), .op(n14679)
         );
  mux2_1 U20327 ( .ip1(\LUT[75][12] ), .ip2(n17544), .s(n17513), .op(n14678)
         );
  mux2_1 U20328 ( .ip1(\LUT[75][11] ), .ip2(n17545), .s(n17513), .op(n14677)
         );
  mux2_1 U20329 ( .ip1(\LUT[75][10] ), .ip2(n17546), .s(n17513), .op(n14676)
         );
  mux2_1 U20330 ( .ip1(\LUT[75][9] ), .ip2(n17547), .s(n17513), .op(n14675) );
  mux2_1 U20331 ( .ip1(\LUT[75][8] ), .ip2(n17548), .s(n17513), .op(n14674) );
  mux2_1 U20332 ( .ip1(\LUT[75][7] ), .ip2(n17549), .s(n17513), .op(n14673) );
  mux2_1 U20333 ( .ip1(\LUT[75][6] ), .ip2(n17551), .s(n17513), .op(n14672) );
  mux2_1 U20334 ( .ip1(\LUT[75][5] ), .ip2(n17552), .s(n17514), .op(n14671) );
  mux2_1 U20335 ( .ip1(\LUT[75][4] ), .ip2(n17553), .s(n17514), .op(n14670) );
  mux2_1 U20336 ( .ip1(\LUT[75][3] ), .ip2(n17554), .s(n17514), .op(n14669) );
  mux2_1 U20337 ( .ip1(\LUT[75][2] ), .ip2(n17555), .s(n17514), .op(n14668) );
  mux2_1 U20338 ( .ip1(\LUT[75][1] ), .ip2(n17556), .s(n17514), .op(n14667) );
  mux2_1 U20339 ( .ip1(\LUT[75][0] ), .ip2(n17558), .s(n17514), .op(n14666) );
  mux2_1 U20340 ( .ip1(\LUT[74][15] ), .ip2(n17541), .s(n17515), .op(n14665)
         );
  mux2_1 U20341 ( .ip1(\LUT[74][14] ), .ip2(n17542), .s(n17515), .op(n14664)
         );
  mux2_1 U20342 ( .ip1(\LUT[74][13] ), .ip2(n17543), .s(n17515), .op(n14663)
         );
  mux2_1 U20343 ( .ip1(\LUT[74][12] ), .ip2(n17544), .s(n17515), .op(n14662)
         );
  mux2_1 U20344 ( .ip1(\LUT[74][11] ), .ip2(n17545), .s(n17515), .op(n14661)
         );
  mux2_1 U20345 ( .ip1(\LUT[74][10] ), .ip2(n17546), .s(n17515), .op(n14660)
         );
  mux2_1 U20346 ( .ip1(\LUT[74][9] ), .ip2(n17547), .s(n17515), .op(n14659) );
  mux2_1 U20347 ( .ip1(\LUT[74][8] ), .ip2(n17548), .s(n17515), .op(n14658) );
  mux2_1 U20348 ( .ip1(\LUT[74][7] ), .ip2(n17549), .s(n17515), .op(n14657) );
  mux2_1 U20349 ( .ip1(\LUT[74][6] ), .ip2(n17551), .s(n17515), .op(n14656) );
  mux2_1 U20350 ( .ip1(\LUT[74][5] ), .ip2(n17552), .s(n17516), .op(n14655) );
  mux2_1 U20351 ( .ip1(\LUT[74][4] ), .ip2(n17553), .s(n17516), .op(n14654) );
  mux2_1 U20352 ( .ip1(\LUT[74][3] ), .ip2(n17554), .s(n17516), .op(n14653) );
  mux2_1 U20353 ( .ip1(\LUT[74][2] ), .ip2(n17555), .s(n17516), .op(n14652) );
  mux2_1 U20354 ( .ip1(\LUT[74][1] ), .ip2(n17556), .s(n17516), .op(n14651) );
  mux2_1 U20355 ( .ip1(\LUT[74][0] ), .ip2(n17558), .s(n17516), .op(n14650) );
  mux2_1 U20356 ( .ip1(\LUT[73][15] ), .ip2(n17541), .s(n17517), .op(n14649)
         );
  mux2_1 U20357 ( .ip1(\LUT[73][14] ), .ip2(n17542), .s(n17517), .op(n14648)
         );
  mux2_1 U20358 ( .ip1(\LUT[73][13] ), .ip2(n17543), .s(n17517), .op(n14647)
         );
  mux2_1 U20359 ( .ip1(\LUT[73][12] ), .ip2(n17544), .s(n17517), .op(n14646)
         );
  mux2_1 U20360 ( .ip1(\LUT[73][11] ), .ip2(n17545), .s(n17517), .op(n14645)
         );
  mux2_1 U20361 ( .ip1(\LUT[73][10] ), .ip2(n17546), .s(n17517), .op(n14644)
         );
  mux2_1 U20362 ( .ip1(\LUT[73][9] ), .ip2(n17547), .s(n17517), .op(n14643) );
  mux2_1 U20363 ( .ip1(\LUT[73][8] ), .ip2(n17548), .s(n17517), .op(n14642) );
  mux2_1 U20364 ( .ip1(\LUT[73][7] ), .ip2(n17549), .s(n17517), .op(n14641) );
  mux2_1 U20365 ( .ip1(\LUT[73][6] ), .ip2(n17551), .s(n17517), .op(n14640) );
  mux2_1 U20366 ( .ip1(\LUT[73][5] ), .ip2(n17552), .s(n17518), .op(n14639) );
  mux2_1 U20367 ( .ip1(\LUT[73][4] ), .ip2(n17553), .s(n17518), .op(n14638) );
  mux2_1 U20368 ( .ip1(\LUT[73][3] ), .ip2(n17554), .s(n17518), .op(n14637) );
  mux2_1 U20369 ( .ip1(\LUT[73][2] ), .ip2(n17555), .s(n17518), .op(n14636) );
  mux2_1 U20370 ( .ip1(\LUT[73][1] ), .ip2(n17556), .s(n17518), .op(n14635) );
  mux2_1 U20371 ( .ip1(\LUT[73][0] ), .ip2(n17558), .s(n17518), .op(n14634) );
  mux2_1 U20372 ( .ip1(\LUT[72][15] ), .ip2(n17541), .s(n17519), .op(n14633)
         );
  mux2_1 U20373 ( .ip1(\LUT[72][14] ), .ip2(n17542), .s(n17519), .op(n14632)
         );
  mux2_1 U20374 ( .ip1(\LUT[72][13] ), .ip2(n17543), .s(n17519), .op(n14631)
         );
  mux2_1 U20375 ( .ip1(\LUT[72][12] ), .ip2(n17544), .s(n17519), .op(n14630)
         );
  mux2_1 U20376 ( .ip1(\LUT[72][11] ), .ip2(n17545), .s(n17519), .op(n14629)
         );
  mux2_1 U20377 ( .ip1(\LUT[72][10] ), .ip2(n17546), .s(n17519), .op(n14628)
         );
  mux2_1 U20378 ( .ip1(\LUT[72][9] ), .ip2(n17547), .s(n17519), .op(n14627) );
  mux2_1 U20379 ( .ip1(\LUT[72][8] ), .ip2(n17548), .s(n17519), .op(n14626) );
  mux2_1 U20380 ( .ip1(\LUT[72][7] ), .ip2(n17549), .s(n17519), .op(n14625) );
  mux2_1 U20381 ( .ip1(\LUT[72][6] ), .ip2(n17551), .s(n17519), .op(n14624) );
  mux2_1 U20382 ( .ip1(\LUT[72][5] ), .ip2(n17552), .s(n17520), .op(n14623) );
  mux2_1 U20383 ( .ip1(\LUT[72][4] ), .ip2(n17553), .s(n17520), .op(n14622) );
  mux2_1 U20384 ( .ip1(\LUT[72][3] ), .ip2(n17554), .s(n17520), .op(n14621) );
  mux2_1 U20385 ( .ip1(\LUT[72][2] ), .ip2(n17555), .s(n17520), .op(n14620) );
  mux2_1 U20386 ( .ip1(\LUT[72][1] ), .ip2(n17556), .s(n17520), .op(n14619) );
  mux2_1 U20387 ( .ip1(\LUT[72][0] ), .ip2(n17558), .s(n17520), .op(n14618) );
  mux2_1 U20388 ( .ip1(\LUT[71][15] ), .ip2(n17541), .s(n17521), .op(n14617)
         );
  mux2_1 U20389 ( .ip1(\LUT[71][14] ), .ip2(n17542), .s(n17521), .op(n14616)
         );
  mux2_1 U20390 ( .ip1(\LUT[71][13] ), .ip2(n17543), .s(n17521), .op(n14615)
         );
  mux2_1 U20391 ( .ip1(\LUT[71][12] ), .ip2(n17544), .s(n17521), .op(n14614)
         );
  mux2_1 U20392 ( .ip1(\LUT[71][11] ), .ip2(n17545), .s(n17521), .op(n14613)
         );
  mux2_1 U20393 ( .ip1(\LUT[71][10] ), .ip2(n17546), .s(n17521), .op(n14612)
         );
  mux2_1 U20394 ( .ip1(\LUT[71][9] ), .ip2(n17547), .s(n17521), .op(n14611) );
  mux2_1 U20395 ( .ip1(\LUT[71][8] ), .ip2(n17548), .s(n17521), .op(n14610) );
  mux2_1 U20396 ( .ip1(\LUT[71][7] ), .ip2(n17549), .s(n17521), .op(n14609) );
  mux2_1 U20397 ( .ip1(\LUT[71][6] ), .ip2(n17551), .s(n17521), .op(n14608) );
  mux2_1 U20398 ( .ip1(\LUT[71][5] ), .ip2(n17552), .s(n17522), .op(n14607) );
  mux2_1 U20399 ( .ip1(\LUT[71][4] ), .ip2(n17553), .s(n17522), .op(n14606) );
  mux2_1 U20400 ( .ip1(\LUT[71][3] ), .ip2(n17554), .s(n17522), .op(n14605) );
  mux2_1 U20401 ( .ip1(\LUT[71][2] ), .ip2(n17555), .s(n17522), .op(n14604) );
  mux2_1 U20402 ( .ip1(\LUT[71][1] ), .ip2(n17556), .s(n17522), .op(n14603) );
  mux2_1 U20403 ( .ip1(\LUT[71][0] ), .ip2(n17558), .s(n17522), .op(n14602) );
  mux2_1 U20404 ( .ip1(\LUT[70][15] ), .ip2(d[15]), .s(n17523), .op(n14601) );
  mux2_1 U20405 ( .ip1(\LUT[70][14] ), .ip2(d[14]), .s(n17523), .op(n14600) );
  mux2_1 U20406 ( .ip1(\LUT[70][13] ), .ip2(d[13]), .s(n17523), .op(n14599) );
  mux2_1 U20407 ( .ip1(\LUT[70][12] ), .ip2(d[12]), .s(n17523), .op(n14598) );
  mux2_1 U20408 ( .ip1(\LUT[70][11] ), .ip2(d[11]), .s(n17523), .op(n14597) );
  mux2_1 U20409 ( .ip1(\LUT[70][10] ), .ip2(d[10]), .s(n17523), .op(n14596) );
  mux2_1 U20410 ( .ip1(\LUT[70][9] ), .ip2(d[9]), .s(n17523), .op(n14595) );
  mux2_1 U20411 ( .ip1(\LUT[70][8] ), .ip2(d[8]), .s(n17523), .op(n14594) );
  mux2_1 U20412 ( .ip1(\LUT[70][7] ), .ip2(d[7]), .s(n17523), .op(n14593) );
  mux2_1 U20413 ( .ip1(\LUT[70][6] ), .ip2(d[6]), .s(n17523), .op(n14592) );
  mux2_1 U20414 ( .ip1(\LUT[70][5] ), .ip2(d[5]), .s(n17524), .op(n14591) );
  mux2_1 U20415 ( .ip1(\LUT[70][4] ), .ip2(d[4]), .s(n17524), .op(n14590) );
  mux2_1 U20416 ( .ip1(\LUT[70][3] ), .ip2(d[3]), .s(n17524), .op(n14589) );
  mux2_1 U20417 ( .ip1(\LUT[70][2] ), .ip2(d[2]), .s(n17524), .op(n14588) );
  mux2_1 U20418 ( .ip1(\LUT[70][1] ), .ip2(d[1]), .s(n17524), .op(n14587) );
  mux2_1 U20419 ( .ip1(\LUT[70][0] ), .ip2(d[0]), .s(n17524), .op(n14586) );
  mux2_1 U20420 ( .ip1(\LUT[69][15] ), .ip2(n17541), .s(n17525), .op(n14585)
         );
  mux2_1 U20421 ( .ip1(\LUT[69][14] ), .ip2(n17542), .s(n17525), .op(n14584)
         );
  mux2_1 U20422 ( .ip1(\LUT[69][13] ), .ip2(n17543), .s(n17525), .op(n14583)
         );
  mux2_1 U20423 ( .ip1(\LUT[69][12] ), .ip2(n17544), .s(n17525), .op(n14582)
         );
  mux2_1 U20424 ( .ip1(\LUT[69][11] ), .ip2(n17545), .s(n17525), .op(n14581)
         );
  mux2_1 U20425 ( .ip1(\LUT[69][10] ), .ip2(n17546), .s(n17525), .op(n14580)
         );
  mux2_1 U20426 ( .ip1(\LUT[69][9] ), .ip2(n17547), .s(n17525), .op(n14579) );
  mux2_1 U20427 ( .ip1(\LUT[69][8] ), .ip2(n17548), .s(n17525), .op(n14578) );
  mux2_1 U20428 ( .ip1(\LUT[69][7] ), .ip2(n17549), .s(n17525), .op(n14577) );
  mux2_1 U20429 ( .ip1(\LUT[69][6] ), .ip2(n17551), .s(n17525), .op(n14576) );
  mux2_1 U20430 ( .ip1(\LUT[69][5] ), .ip2(n17552), .s(n17526), .op(n14575) );
  mux2_1 U20431 ( .ip1(\LUT[69][4] ), .ip2(n17553), .s(n17526), .op(n14574) );
  mux2_1 U20432 ( .ip1(\LUT[69][3] ), .ip2(n17554), .s(n17526), .op(n14573) );
  mux2_1 U20433 ( .ip1(\LUT[69][2] ), .ip2(n17555), .s(n17526), .op(n14572) );
  mux2_1 U20434 ( .ip1(\LUT[69][1] ), .ip2(n17556), .s(n17526), .op(n14571) );
  mux2_1 U20435 ( .ip1(\LUT[69][0] ), .ip2(n17558), .s(n17526), .op(n14570) );
  mux2_1 U20436 ( .ip1(\LUT[68][15] ), .ip2(d[15]), .s(n17527), .op(n14569) );
  mux2_1 U20437 ( .ip1(\LUT[68][14] ), .ip2(d[14]), .s(n17527), .op(n14568) );
  mux2_1 U20438 ( .ip1(\LUT[68][13] ), .ip2(d[13]), .s(n17527), .op(n14567) );
  mux2_1 U20439 ( .ip1(\LUT[68][12] ), .ip2(d[12]), .s(n17527), .op(n14566) );
  mux2_1 U20440 ( .ip1(\LUT[68][11] ), .ip2(d[11]), .s(n17527), .op(n14565) );
  mux2_1 U20441 ( .ip1(\LUT[68][10] ), .ip2(d[10]), .s(n17527), .op(n14564) );
  mux2_1 U20442 ( .ip1(\LUT[68][9] ), .ip2(d[9]), .s(n17527), .op(n14563) );
  mux2_1 U20443 ( .ip1(\LUT[68][8] ), .ip2(d[8]), .s(n17527), .op(n14562) );
  mux2_1 U20444 ( .ip1(\LUT[68][7] ), .ip2(d[7]), .s(n17527), .op(n14561) );
  mux2_1 U20445 ( .ip1(\LUT[68][6] ), .ip2(d[6]), .s(n17527), .op(n14560) );
  mux2_1 U20446 ( .ip1(\LUT[68][5] ), .ip2(d[5]), .s(n17528), .op(n14559) );
  mux2_1 U20447 ( .ip1(\LUT[68][4] ), .ip2(d[4]), .s(n17528), .op(n14558) );
  mux2_1 U20448 ( .ip1(\LUT[68][3] ), .ip2(d[3]), .s(n17528), .op(n14557) );
  mux2_1 U20449 ( .ip1(\LUT[68][2] ), .ip2(d[2]), .s(n17528), .op(n14556) );
  mux2_1 U20450 ( .ip1(\LUT[68][1] ), .ip2(d[1]), .s(n17528), .op(n14555) );
  mux2_1 U20451 ( .ip1(\LUT[68][0] ), .ip2(d[0]), .s(n17528), .op(n14554) );
  mux2_1 U20452 ( .ip1(\LUT[67][15] ), .ip2(n17541), .s(n17529), .op(n14553)
         );
  mux2_1 U20453 ( .ip1(\LUT[67][14] ), .ip2(n17542), .s(n17529), .op(n14552)
         );
  mux2_1 U20454 ( .ip1(\LUT[67][13] ), .ip2(n17543), .s(n17529), .op(n14551)
         );
  mux2_1 U20455 ( .ip1(\LUT[67][12] ), .ip2(n17544), .s(n17529), .op(n14550)
         );
  mux2_1 U20456 ( .ip1(\LUT[67][11] ), .ip2(n17545), .s(n17529), .op(n14549)
         );
  mux2_1 U20457 ( .ip1(\LUT[67][10] ), .ip2(n17546), .s(n17529), .op(n14548)
         );
  mux2_1 U20458 ( .ip1(\LUT[67][9] ), .ip2(n17547), .s(n17529), .op(n14547) );
  mux2_1 U20459 ( .ip1(\LUT[67][8] ), .ip2(n17548), .s(n17529), .op(n14546) );
  mux2_1 U20460 ( .ip1(\LUT[67][7] ), .ip2(n17549), .s(n17529), .op(n14545) );
  mux2_1 U20461 ( .ip1(\LUT[67][6] ), .ip2(n17551), .s(n17529), .op(n14544) );
  mux2_1 U20462 ( .ip1(\LUT[67][5] ), .ip2(n17552), .s(n17530), .op(n14543) );
  mux2_1 U20463 ( .ip1(\LUT[67][4] ), .ip2(n17553), .s(n17530), .op(n14542) );
  mux2_1 U20464 ( .ip1(\LUT[67][3] ), .ip2(n17554), .s(n17530), .op(n14541) );
  mux2_1 U20465 ( .ip1(\LUT[67][2] ), .ip2(n17555), .s(n17530), .op(n14540) );
  mux2_1 U20466 ( .ip1(\LUT[67][1] ), .ip2(n17556), .s(n17530), .op(n14539) );
  mux2_1 U20467 ( .ip1(\LUT[67][0] ), .ip2(n17558), .s(n17530), .op(n14538) );
  mux2_1 U20468 ( .ip1(\LUT[66][15] ), .ip2(d[15]), .s(n17531), .op(n14537) );
  mux2_1 U20469 ( .ip1(\LUT[66][14] ), .ip2(d[14]), .s(n17531), .op(n14536) );
  mux2_1 U20470 ( .ip1(\LUT[66][13] ), .ip2(d[13]), .s(n17531), .op(n14535) );
  mux2_1 U20471 ( .ip1(\LUT[66][12] ), .ip2(d[12]), .s(n17531), .op(n14534) );
  mux2_1 U20472 ( .ip1(\LUT[66][11] ), .ip2(d[11]), .s(n17531), .op(n14533) );
  mux2_1 U20473 ( .ip1(\LUT[66][10] ), .ip2(d[10]), .s(n17531), .op(n14532) );
  mux2_1 U20474 ( .ip1(\LUT[66][9] ), .ip2(d[9]), .s(n17531), .op(n14531) );
  mux2_1 U20475 ( .ip1(\LUT[66][8] ), .ip2(d[8]), .s(n17531), .op(n14530) );
  mux2_1 U20476 ( .ip1(\LUT[66][7] ), .ip2(d[7]), .s(n17531), .op(n14529) );
  mux2_1 U20477 ( .ip1(\LUT[66][6] ), .ip2(d[6]), .s(n17531), .op(n14528) );
  mux2_1 U20478 ( .ip1(\LUT[66][5] ), .ip2(d[5]), .s(n17532), .op(n14527) );
  mux2_1 U20479 ( .ip1(\LUT[66][4] ), .ip2(d[4]), .s(n17532), .op(n14526) );
  mux2_1 U20480 ( .ip1(\LUT[66][3] ), .ip2(d[3]), .s(n17532), .op(n14525) );
  mux2_1 U20481 ( .ip1(\LUT[66][2] ), .ip2(d[2]), .s(n17532), .op(n14524) );
  mux2_1 U20482 ( .ip1(\LUT[66][1] ), .ip2(d[1]), .s(n17532), .op(n14523) );
  mux2_1 U20483 ( .ip1(\LUT[66][0] ), .ip2(d[0]), .s(n17532), .op(n14522) );
  mux2_1 U20484 ( .ip1(\LUT[65][15] ), .ip2(n17541), .s(n17533), .op(n14521)
         );
  mux2_1 U20485 ( .ip1(\LUT[65][14] ), .ip2(n17542), .s(n17533), .op(n14520)
         );
  mux2_1 U20486 ( .ip1(\LUT[65][13] ), .ip2(n17543), .s(n17533), .op(n14519)
         );
  mux2_1 U20487 ( .ip1(\LUT[65][12] ), .ip2(n17544), .s(n17533), .op(n14518)
         );
  mux2_1 U20488 ( .ip1(\LUT[65][11] ), .ip2(n17545), .s(n17533), .op(n14517)
         );
  mux2_1 U20489 ( .ip1(\LUT[65][10] ), .ip2(n17546), .s(n17533), .op(n14516)
         );
  mux2_1 U20490 ( .ip1(\LUT[65][9] ), .ip2(n17547), .s(n17533), .op(n14515) );
  mux2_1 U20491 ( .ip1(\LUT[65][8] ), .ip2(n17548), .s(n17533), .op(n14514) );
  mux2_1 U20492 ( .ip1(\LUT[65][7] ), .ip2(n17549), .s(n17533), .op(n14513) );
  mux2_1 U20493 ( .ip1(\LUT[65][6] ), .ip2(n17551), .s(n17533), .op(n14512) );
  mux2_1 U20494 ( .ip1(\LUT[65][5] ), .ip2(n17552), .s(n17534), .op(n14511) );
  mux2_1 U20495 ( .ip1(\LUT[65][4] ), .ip2(n17553), .s(n17534), .op(n14510) );
  mux2_1 U20496 ( .ip1(\LUT[65][3] ), .ip2(n17554), .s(n17534), .op(n14509) );
  mux2_1 U20497 ( .ip1(\LUT[65][2] ), .ip2(n17555), .s(n17534), .op(n14508) );
  mux2_1 U20498 ( .ip1(\LUT[65][1] ), .ip2(n17556), .s(n17534), .op(n14507) );
  mux2_1 U20499 ( .ip1(\LUT[65][0] ), .ip2(n17558), .s(n17534), .op(n14506) );
  mux2_1 U20500 ( .ip1(\LUT[64][15] ), .ip2(d[15]), .s(n17535), .op(n14505) );
  mux2_1 U20501 ( .ip1(\LUT[64][14] ), .ip2(d[14]), .s(n17535), .op(n14504) );
  mux2_1 U20502 ( .ip1(\LUT[64][13] ), .ip2(d[13]), .s(n17535), .op(n14503) );
  mux2_1 U20503 ( .ip1(\LUT[64][12] ), .ip2(d[12]), .s(n17535), .op(n14502) );
  mux2_1 U20504 ( .ip1(\LUT[64][11] ), .ip2(d[11]), .s(n17535), .op(n14501) );
  mux2_1 U20505 ( .ip1(\LUT[64][10] ), .ip2(d[10]), .s(n17535), .op(n14500) );
  mux2_1 U20506 ( .ip1(\LUT[64][9] ), .ip2(d[9]), .s(n17535), .op(n14499) );
  mux2_1 U20507 ( .ip1(\LUT[64][8] ), .ip2(d[8]), .s(n17535), .op(n14498) );
  mux2_1 U20508 ( .ip1(\LUT[64][7] ), .ip2(d[7]), .s(n17535), .op(n14497) );
  mux2_1 U20509 ( .ip1(\LUT[64][6] ), .ip2(d[6]), .s(n17535), .op(n14496) );
  mux2_1 U20510 ( .ip1(\LUT[64][5] ), .ip2(d[5]), .s(n17536), .op(n14495) );
  mux2_1 U20511 ( .ip1(\LUT[64][4] ), .ip2(d[4]), .s(n17536), .op(n14494) );
  mux2_1 U20512 ( .ip1(\LUT[64][3] ), .ip2(d[3]), .s(n17536), .op(n14493) );
  mux2_1 U20513 ( .ip1(\LUT[64][2] ), .ip2(d[2]), .s(n17536), .op(n14492) );
  mux2_1 U20514 ( .ip1(\LUT[64][1] ), .ip2(d[1]), .s(n17536), .op(n14491) );
  mux2_1 U20515 ( .ip1(\LUT[64][0] ), .ip2(d[0]), .s(n17536), .op(n14490) );
  mux2_1 U20516 ( .ip1(\LUT[63][15] ), .ip2(n17541), .s(n17537), .op(n14489)
         );
  mux2_1 U20517 ( .ip1(\LUT[63][14] ), .ip2(n17542), .s(n17537), .op(n14488)
         );
  mux2_1 U20518 ( .ip1(\LUT[63][13] ), .ip2(n17543), .s(n17537), .op(n14487)
         );
  mux2_1 U20519 ( .ip1(\LUT[63][12] ), .ip2(n17544), .s(n17537), .op(n14486)
         );
  mux2_1 U20520 ( .ip1(\LUT[63][11] ), .ip2(n17545), .s(n17537), .op(n14485)
         );
  mux2_1 U20521 ( .ip1(\LUT[63][10] ), .ip2(n17546), .s(n17537), .op(n14484)
         );
  mux2_1 U20522 ( .ip1(\LUT[63][9] ), .ip2(n17547), .s(n17537), .op(n14483) );
  mux2_1 U20523 ( .ip1(\LUT[63][8] ), .ip2(n17548), .s(n17537), .op(n14482) );
  mux2_1 U20524 ( .ip1(\LUT[63][7] ), .ip2(n17549), .s(n17537), .op(n14481) );
  mux2_1 U20525 ( .ip1(\LUT[63][6] ), .ip2(n17551), .s(n17537), .op(n14480) );
  mux2_1 U20526 ( .ip1(\LUT[63][5] ), .ip2(n17552), .s(n17538), .op(n14479) );
  mux2_1 U20527 ( .ip1(\LUT[63][4] ), .ip2(n17553), .s(n17538), .op(n14478) );
  mux2_1 U20528 ( .ip1(\LUT[63][3] ), .ip2(n17554), .s(n17538), .op(n14477) );
  mux2_1 U20529 ( .ip1(\LUT[63][2] ), .ip2(n17555), .s(n17538), .op(n14476) );
  mux2_1 U20530 ( .ip1(\LUT[63][1] ), .ip2(n17556), .s(n17538), .op(n14475) );
  mux2_1 U20531 ( .ip1(\LUT[63][0] ), .ip2(n17558), .s(n17538), .op(n14474) );
  mux2_1 U20532 ( .ip1(\LUT[62][15] ), .ip2(d[15]), .s(n17539), .op(n14473) );
  mux2_1 U20533 ( .ip1(\LUT[62][14] ), .ip2(d[14]), .s(n17539), .op(n14472) );
  mux2_1 U20534 ( .ip1(\LUT[62][13] ), .ip2(d[13]), .s(n17539), .op(n14471) );
  mux2_1 U20535 ( .ip1(\LUT[62][12] ), .ip2(d[12]), .s(n17539), .op(n14470) );
  mux2_1 U20536 ( .ip1(\LUT[62][11] ), .ip2(d[11]), .s(n17539), .op(n14469) );
  mux2_1 U20537 ( .ip1(\LUT[62][10] ), .ip2(d[10]), .s(n17539), .op(n14468) );
  mux2_1 U20538 ( .ip1(\LUT[62][9] ), .ip2(d[9]), .s(n17539), .op(n14467) );
  mux2_1 U20539 ( .ip1(\LUT[62][8] ), .ip2(d[8]), .s(n17539), .op(n14466) );
  mux2_1 U20540 ( .ip1(\LUT[62][7] ), .ip2(d[7]), .s(n17539), .op(n14465) );
  mux2_1 U20541 ( .ip1(\LUT[62][6] ), .ip2(d[6]), .s(n17539), .op(n14464) );
  mux2_1 U20542 ( .ip1(\LUT[62][5] ), .ip2(d[5]), .s(n17540), .op(n14463) );
  mux2_1 U20543 ( .ip1(\LUT[62][4] ), .ip2(d[4]), .s(n17540), .op(n14462) );
  mux2_1 U20544 ( .ip1(\LUT[62][3] ), .ip2(d[3]), .s(n17540), .op(n14461) );
  mux2_1 U20545 ( .ip1(\LUT[62][2] ), .ip2(d[2]), .s(n17540), .op(n14460) );
  mux2_1 U20546 ( .ip1(\LUT[62][1] ), .ip2(d[1]), .s(n17540), .op(n14459) );
  mux2_1 U20547 ( .ip1(\LUT[62][0] ), .ip2(d[0]), .s(n17540), .op(n14458) );
  mux2_1 U20548 ( .ip1(\LUT[61][15] ), .ip2(n17541), .s(n17550), .op(n14457)
         );
  mux2_1 U20549 ( .ip1(\LUT[61][14] ), .ip2(n17542), .s(n17550), .op(n14456)
         );
  mux2_1 U20550 ( .ip1(\LUT[61][13] ), .ip2(n17543), .s(n17550), .op(n14455)
         );
  mux2_1 U20551 ( .ip1(\LUT[61][12] ), .ip2(n17544), .s(n17550), .op(n14454)
         );
  mux2_1 U20552 ( .ip1(\LUT[61][11] ), .ip2(n17545), .s(n17550), .op(n14453)
         );
  mux2_1 U20553 ( .ip1(\LUT[61][10] ), .ip2(n17546), .s(n17550), .op(n14452)
         );
  mux2_1 U20554 ( .ip1(\LUT[61][9] ), .ip2(n17547), .s(n17550), .op(n14451) );
  mux2_1 U20555 ( .ip1(\LUT[61][8] ), .ip2(n17548), .s(n17550), .op(n14450) );
  mux2_1 U20556 ( .ip1(\LUT[61][7] ), .ip2(n17549), .s(n17550), .op(n14449) );
  mux2_1 U20557 ( .ip1(\LUT[61][6] ), .ip2(n17551), .s(n17550), .op(n14448) );
  mux2_1 U20558 ( .ip1(\LUT[61][5] ), .ip2(n17552), .s(n17557), .op(n14447) );
  mux2_1 U20559 ( .ip1(\LUT[61][4] ), .ip2(n17553), .s(n17557), .op(n14446) );
  mux2_1 U20560 ( .ip1(\LUT[61][3] ), .ip2(n17554), .s(n17557), .op(n14445) );
  mux2_1 U20561 ( .ip1(\LUT[61][2] ), .ip2(n17555), .s(n17557), .op(n14444) );
  mux2_1 U20562 ( .ip1(\LUT[61][1] ), .ip2(n17556), .s(n17557), .op(n14443) );
  mux2_1 U20563 ( .ip1(\LUT[61][0] ), .ip2(n17558), .s(n17557), .op(n14442) );
  buf_1 U20564 ( .ip(d[15]), .op(n17629) );
  mux2_1 U20565 ( .ip1(\LUT[60][15] ), .ip2(n17629), .s(n17559), .op(n14441)
         );
  buf_1 U20566 ( .ip(d[14]), .op(n17630) );
  mux2_1 U20567 ( .ip1(\LUT[60][14] ), .ip2(n17630), .s(n17559), .op(n14440)
         );
  buf_1 U20568 ( .ip(d[13]), .op(n17631) );
  mux2_1 U20569 ( .ip1(\LUT[60][13] ), .ip2(n17631), .s(n17559), .op(n14439)
         );
  buf_1 U20570 ( .ip(d[12]), .op(n17632) );
  mux2_1 U20571 ( .ip1(\LUT[60][12] ), .ip2(n17632), .s(n17559), .op(n14438)
         );
  buf_1 U20572 ( .ip(d[11]), .op(n17633) );
  mux2_1 U20573 ( .ip1(\LUT[60][11] ), .ip2(n17633), .s(n17559), .op(n14437)
         );
  buf_1 U20574 ( .ip(d[10]), .op(n17634) );
  mux2_1 U20575 ( .ip1(\LUT[60][10] ), .ip2(n17634), .s(n17559), .op(n14436)
         );
  buf_1 U20576 ( .ip(d[9]), .op(n17635) );
  mux2_1 U20577 ( .ip1(\LUT[60][9] ), .ip2(n17635), .s(n17559), .op(n14435) );
  buf_1 U20578 ( .ip(d[8]), .op(n17636) );
  mux2_1 U20579 ( .ip1(\LUT[60][8] ), .ip2(n17636), .s(n17559), .op(n14434) );
  buf_1 U20580 ( .ip(d[7]), .op(n17637) );
  mux2_1 U20581 ( .ip1(\LUT[60][7] ), .ip2(n17637), .s(n17559), .op(n14433) );
  buf_1 U20582 ( .ip(d[6]), .op(n17639) );
  mux2_1 U20583 ( .ip1(\LUT[60][6] ), .ip2(n17639), .s(n17559), .op(n14432) );
  buf_1 U20584 ( .ip(d[5]), .op(n17640) );
  mux2_1 U20585 ( .ip1(\LUT[60][5] ), .ip2(n17640), .s(n17560), .op(n14431) );
  buf_1 U20586 ( .ip(d[4]), .op(n17641) );
  mux2_1 U20587 ( .ip1(\LUT[60][4] ), .ip2(n17641), .s(n17560), .op(n14430) );
  buf_1 U20588 ( .ip(d[3]), .op(n17642) );
  mux2_1 U20589 ( .ip1(\LUT[60][3] ), .ip2(n17642), .s(n17560), .op(n14429) );
  buf_1 U20590 ( .ip(d[2]), .op(n17643) );
  mux2_1 U20591 ( .ip1(\LUT[60][2] ), .ip2(n17643), .s(n17560), .op(n14428) );
  buf_1 U20592 ( .ip(d[1]), .op(n17644) );
  mux2_1 U20593 ( .ip1(\LUT[60][1] ), .ip2(n17644), .s(n17560), .op(n14427) );
  buf_1 U20594 ( .ip(d[0]), .op(n17646) );
  mux2_1 U20595 ( .ip1(\LUT[60][0] ), .ip2(n17646), .s(n17560), .op(n14426) );
  mux2_1 U20596 ( .ip1(\LUT[59][15] ), .ip2(n17629), .s(n17561), .op(n14425)
         );
  mux2_1 U20597 ( .ip1(\LUT[59][14] ), .ip2(n17630), .s(n17561), .op(n14424)
         );
  mux2_1 U20598 ( .ip1(\LUT[59][13] ), .ip2(n17631), .s(n17561), .op(n14423)
         );
  mux2_1 U20599 ( .ip1(\LUT[59][12] ), .ip2(n17632), .s(n17561), .op(n14422)
         );
  mux2_1 U20600 ( .ip1(\LUT[59][11] ), .ip2(n17633), .s(n17561), .op(n14421)
         );
  mux2_1 U20601 ( .ip1(\LUT[59][10] ), .ip2(n17634), .s(n17561), .op(n14420)
         );
  mux2_1 U20602 ( .ip1(\LUT[59][9] ), .ip2(n17635), .s(n17561), .op(n14419) );
  mux2_1 U20603 ( .ip1(\LUT[59][8] ), .ip2(n17636), .s(n17561), .op(n14418) );
  mux2_1 U20604 ( .ip1(\LUT[59][7] ), .ip2(n17637), .s(n17561), .op(n14417) );
  mux2_1 U20605 ( .ip1(\LUT[59][6] ), .ip2(n17639), .s(n17561), .op(n14416) );
  mux2_1 U20606 ( .ip1(\LUT[59][5] ), .ip2(n17640), .s(n17562), .op(n14415) );
  mux2_1 U20607 ( .ip1(\LUT[59][4] ), .ip2(n17641), .s(n17562), .op(n14414) );
  mux2_1 U20608 ( .ip1(\LUT[59][3] ), .ip2(n17642), .s(n17562), .op(n14413) );
  mux2_1 U20609 ( .ip1(\LUT[59][2] ), .ip2(n17643), .s(n17562), .op(n14412) );
  mux2_1 U20610 ( .ip1(\LUT[59][1] ), .ip2(n17644), .s(n17562), .op(n14411) );
  mux2_1 U20611 ( .ip1(\LUT[59][0] ), .ip2(n17646), .s(n17562), .op(n14410) );
  mux2_1 U20612 ( .ip1(\LUT[58][15] ), .ip2(n17629), .s(n17563), .op(n14409)
         );
  mux2_1 U20613 ( .ip1(\LUT[58][14] ), .ip2(n17630), .s(n17563), .op(n14408)
         );
  mux2_1 U20614 ( .ip1(\LUT[58][13] ), .ip2(n17631), .s(n17563), .op(n14407)
         );
  mux2_1 U20615 ( .ip1(\LUT[58][12] ), .ip2(n17632), .s(n17563), .op(n14406)
         );
  mux2_1 U20616 ( .ip1(\LUT[58][11] ), .ip2(n17633), .s(n17563), .op(n14405)
         );
  mux2_1 U20617 ( .ip1(\LUT[58][10] ), .ip2(n17634), .s(n17563), .op(n14404)
         );
  mux2_1 U20618 ( .ip1(\LUT[58][9] ), .ip2(n17635), .s(n17563), .op(n14403) );
  mux2_1 U20619 ( .ip1(\LUT[58][8] ), .ip2(n17636), .s(n17563), .op(n14402) );
  mux2_1 U20620 ( .ip1(\LUT[58][7] ), .ip2(n17637), .s(n17563), .op(n14401) );
  mux2_1 U20621 ( .ip1(\LUT[58][6] ), .ip2(n17639), .s(n17563), .op(n14400) );
  mux2_1 U20622 ( .ip1(\LUT[58][5] ), .ip2(n17640), .s(n17564), .op(n14399) );
  mux2_1 U20623 ( .ip1(\LUT[58][4] ), .ip2(n17641), .s(n17564), .op(n14398) );
  mux2_1 U20624 ( .ip1(\LUT[58][3] ), .ip2(n17642), .s(n17564), .op(n14397) );
  mux2_1 U20625 ( .ip1(\LUT[58][2] ), .ip2(n17643), .s(n17564), .op(n14396) );
  mux2_1 U20626 ( .ip1(\LUT[58][1] ), .ip2(n17644), .s(n17564), .op(n14395) );
  mux2_1 U20627 ( .ip1(\LUT[58][0] ), .ip2(n17646), .s(n17564), .op(n14394) );
  mux2_1 U20628 ( .ip1(\LUT[57][15] ), .ip2(n17629), .s(n17565), .op(n14393)
         );
  mux2_1 U20629 ( .ip1(\LUT[57][14] ), .ip2(n17630), .s(n17565), .op(n14392)
         );
  mux2_1 U20630 ( .ip1(\LUT[57][13] ), .ip2(n17631), .s(n17565), .op(n14391)
         );
  mux2_1 U20631 ( .ip1(\LUT[57][12] ), .ip2(n17632), .s(n17565), .op(n14390)
         );
  mux2_1 U20632 ( .ip1(\LUT[57][11] ), .ip2(n17633), .s(n17565), .op(n14389)
         );
  mux2_1 U20633 ( .ip1(\LUT[57][10] ), .ip2(n17634), .s(n17565), .op(n14388)
         );
  mux2_1 U20634 ( .ip1(\LUT[57][9] ), .ip2(n17635), .s(n17565), .op(n14387) );
  mux2_1 U20635 ( .ip1(\LUT[57][8] ), .ip2(n17636), .s(n17565), .op(n14386) );
  mux2_1 U20636 ( .ip1(\LUT[57][7] ), .ip2(n17637), .s(n17565), .op(n14385) );
  mux2_1 U20637 ( .ip1(\LUT[57][6] ), .ip2(n17639), .s(n17565), .op(n14384) );
  mux2_1 U20638 ( .ip1(\LUT[57][5] ), .ip2(n17640), .s(n17566), .op(n14383) );
  mux2_1 U20639 ( .ip1(\LUT[57][4] ), .ip2(n17641), .s(n17566), .op(n14382) );
  mux2_1 U20640 ( .ip1(\LUT[57][3] ), .ip2(n17642), .s(n17566), .op(n14381) );
  mux2_1 U20641 ( .ip1(\LUT[57][2] ), .ip2(n17643), .s(n17566), .op(n14380) );
  mux2_1 U20642 ( .ip1(\LUT[57][1] ), .ip2(n17644), .s(n17566), .op(n14379) );
  mux2_1 U20643 ( .ip1(\LUT[57][0] ), .ip2(n17646), .s(n17566), .op(n14378) );
  mux2_1 U20644 ( .ip1(\LUT[56][15] ), .ip2(n17629), .s(n17567), .op(n14377)
         );
  mux2_1 U20645 ( .ip1(\LUT[56][14] ), .ip2(n17630), .s(n17567), .op(n14376)
         );
  mux2_1 U20646 ( .ip1(\LUT[56][13] ), .ip2(n17631), .s(n17567), .op(n14375)
         );
  mux2_1 U20647 ( .ip1(\LUT[56][12] ), .ip2(n17632), .s(n17567), .op(n14374)
         );
  mux2_1 U20648 ( .ip1(\LUT[56][11] ), .ip2(n17633), .s(n17567), .op(n14373)
         );
  mux2_1 U20649 ( .ip1(\LUT[56][10] ), .ip2(n17634), .s(n17567), .op(n14372)
         );
  mux2_1 U20650 ( .ip1(\LUT[56][9] ), .ip2(n17635), .s(n17567), .op(n14371) );
  mux2_1 U20651 ( .ip1(\LUT[56][8] ), .ip2(n17636), .s(n17567), .op(n14370) );
  mux2_1 U20652 ( .ip1(\LUT[56][7] ), .ip2(n17637), .s(n17567), .op(n14369) );
  mux2_1 U20653 ( .ip1(\LUT[56][6] ), .ip2(n17639), .s(n17567), .op(n14368) );
  mux2_1 U20654 ( .ip1(\LUT[56][5] ), .ip2(n17640), .s(n17568), .op(n14367) );
  mux2_1 U20655 ( .ip1(\LUT[56][4] ), .ip2(n17641), .s(n17568), .op(n14366) );
  mux2_1 U20656 ( .ip1(\LUT[56][3] ), .ip2(n17642), .s(n17568), .op(n14365) );
  mux2_1 U20657 ( .ip1(\LUT[56][2] ), .ip2(n17643), .s(n17568), .op(n14364) );
  mux2_1 U20658 ( .ip1(\LUT[56][1] ), .ip2(n17644), .s(n17568), .op(n14363) );
  mux2_1 U20659 ( .ip1(\LUT[56][0] ), .ip2(n17646), .s(n17568), .op(n14362) );
  mux2_1 U20660 ( .ip1(\LUT[55][15] ), .ip2(n17629), .s(n17569), .op(n14361)
         );
  mux2_1 U20661 ( .ip1(\LUT[55][14] ), .ip2(n17630), .s(n17569), .op(n14360)
         );
  mux2_1 U20662 ( .ip1(\LUT[55][13] ), .ip2(n17631), .s(n17569), .op(n14359)
         );
  mux2_1 U20663 ( .ip1(\LUT[55][12] ), .ip2(n17632), .s(n17569), .op(n14358)
         );
  mux2_1 U20664 ( .ip1(\LUT[55][11] ), .ip2(n17633), .s(n17569), .op(n14357)
         );
  mux2_1 U20665 ( .ip1(\LUT[55][10] ), .ip2(n17634), .s(n17569), .op(n14356)
         );
  mux2_1 U20666 ( .ip1(\LUT[55][9] ), .ip2(n17635), .s(n17569), .op(n14355) );
  mux2_1 U20667 ( .ip1(\LUT[55][8] ), .ip2(n17636), .s(n17569), .op(n14354) );
  mux2_1 U20668 ( .ip1(\LUT[55][7] ), .ip2(n17637), .s(n17569), .op(n14353) );
  mux2_1 U20669 ( .ip1(\LUT[55][6] ), .ip2(n17639), .s(n17569), .op(n14352) );
  mux2_1 U20670 ( .ip1(\LUT[55][5] ), .ip2(n17640), .s(n17570), .op(n14351) );
  mux2_1 U20671 ( .ip1(\LUT[55][4] ), .ip2(n17641), .s(n17570), .op(n14350) );
  mux2_1 U20672 ( .ip1(\LUT[55][3] ), .ip2(n17642), .s(n17570), .op(n14349) );
  mux2_1 U20673 ( .ip1(\LUT[55][2] ), .ip2(n17643), .s(n17570), .op(n14348) );
  mux2_1 U20674 ( .ip1(\LUT[55][1] ), .ip2(n17644), .s(n17570), .op(n14347) );
  mux2_1 U20675 ( .ip1(\LUT[55][0] ), .ip2(n17646), .s(n17570), .op(n14346) );
  mux2_1 U20676 ( .ip1(\LUT[54][15] ), .ip2(n17629), .s(n17571), .op(n14345)
         );
  mux2_1 U20677 ( .ip1(\LUT[54][14] ), .ip2(n17630), .s(n17571), .op(n14344)
         );
  mux2_1 U20678 ( .ip1(\LUT[54][13] ), .ip2(n17631), .s(n17571), .op(n14343)
         );
  mux2_1 U20679 ( .ip1(\LUT[54][12] ), .ip2(n17632), .s(n17571), .op(n14342)
         );
  mux2_1 U20680 ( .ip1(\LUT[54][11] ), .ip2(n17633), .s(n17571), .op(n14341)
         );
  mux2_1 U20681 ( .ip1(\LUT[54][10] ), .ip2(n17634), .s(n17571), .op(n14340)
         );
  mux2_1 U20682 ( .ip1(\LUT[54][9] ), .ip2(n17635), .s(n17571), .op(n14339) );
  mux2_1 U20683 ( .ip1(\LUT[54][8] ), .ip2(n17636), .s(n17571), .op(n14338) );
  mux2_1 U20684 ( .ip1(\LUT[54][7] ), .ip2(n17637), .s(n17571), .op(n14337) );
  mux2_1 U20685 ( .ip1(\LUT[54][6] ), .ip2(n17639), .s(n17571), .op(n14336) );
  mux2_1 U20686 ( .ip1(\LUT[54][5] ), .ip2(n17640), .s(n17572), .op(n14335) );
  mux2_1 U20687 ( .ip1(\LUT[54][4] ), .ip2(n17641), .s(n17572), .op(n14334) );
  mux2_1 U20688 ( .ip1(\LUT[54][3] ), .ip2(n17642), .s(n17572), .op(n14333) );
  mux2_1 U20689 ( .ip1(\LUT[54][2] ), .ip2(n17643), .s(n17572), .op(n14332) );
  mux2_1 U20690 ( .ip1(\LUT[54][1] ), .ip2(n17644), .s(n17572), .op(n14331) );
  mux2_1 U20691 ( .ip1(\LUT[54][0] ), .ip2(n17646), .s(n17572), .op(n14330) );
  mux2_1 U20692 ( .ip1(\LUT[53][15] ), .ip2(n17629), .s(n17573), .op(n14329)
         );
  mux2_1 U20693 ( .ip1(\LUT[53][14] ), .ip2(n17630), .s(n17573), .op(n14328)
         );
  mux2_1 U20694 ( .ip1(\LUT[53][13] ), .ip2(n17631), .s(n17573), .op(n14327)
         );
  mux2_1 U20695 ( .ip1(\LUT[53][12] ), .ip2(n17632), .s(n17573), .op(n14326)
         );
  mux2_1 U20696 ( .ip1(\LUT[53][11] ), .ip2(n17633), .s(n17573), .op(n14325)
         );
  mux2_1 U20697 ( .ip1(\LUT[53][10] ), .ip2(n17634), .s(n17573), .op(n14324)
         );
  mux2_1 U20698 ( .ip1(\LUT[53][9] ), .ip2(n17635), .s(n17573), .op(n14323) );
  mux2_1 U20699 ( .ip1(\LUT[53][8] ), .ip2(n17636), .s(n17573), .op(n14322) );
  mux2_1 U20700 ( .ip1(\LUT[53][7] ), .ip2(n17637), .s(n17573), .op(n14321) );
  mux2_1 U20701 ( .ip1(\LUT[53][6] ), .ip2(n17639), .s(n17573), .op(n14320) );
  mux2_1 U20702 ( .ip1(\LUT[53][5] ), .ip2(n17640), .s(n17574), .op(n14319) );
  mux2_1 U20703 ( .ip1(\LUT[53][4] ), .ip2(n17641), .s(n17574), .op(n14318) );
  mux2_1 U20704 ( .ip1(\LUT[53][3] ), .ip2(n17642), .s(n17574), .op(n14317) );
  mux2_1 U20705 ( .ip1(\LUT[53][2] ), .ip2(n17643), .s(n17574), .op(n14316) );
  mux2_1 U20706 ( .ip1(\LUT[53][1] ), .ip2(n17644), .s(n17574), .op(n14315) );
  mux2_1 U20707 ( .ip1(\LUT[53][0] ), .ip2(n17646), .s(n17574), .op(n14314) );
  mux2_1 U20708 ( .ip1(\LUT[52][15] ), .ip2(n17629), .s(n17575), .op(n14313)
         );
  mux2_1 U20709 ( .ip1(\LUT[52][14] ), .ip2(n17630), .s(n17575), .op(n14312)
         );
  mux2_1 U20710 ( .ip1(\LUT[52][13] ), .ip2(n17631), .s(n17575), .op(n14311)
         );
  mux2_1 U20711 ( .ip1(\LUT[52][12] ), .ip2(n17632), .s(n17575), .op(n14310)
         );
  mux2_1 U20712 ( .ip1(\LUT[52][11] ), .ip2(n17633), .s(n17575), .op(n14309)
         );
  mux2_1 U20713 ( .ip1(\LUT[52][10] ), .ip2(n17634), .s(n17575), .op(n14308)
         );
  mux2_1 U20714 ( .ip1(\LUT[52][9] ), .ip2(n17635), .s(n17575), .op(n14307) );
  mux2_1 U20715 ( .ip1(\LUT[52][8] ), .ip2(n17636), .s(n17575), .op(n14306) );
  mux2_1 U20716 ( .ip1(\LUT[52][7] ), .ip2(n17637), .s(n17575), .op(n14305) );
  mux2_1 U20717 ( .ip1(\LUT[52][6] ), .ip2(n17639), .s(n17575), .op(n14304) );
  mux2_1 U20718 ( .ip1(\LUT[52][5] ), .ip2(n17640), .s(n17576), .op(n14303) );
  mux2_1 U20719 ( .ip1(\LUT[52][4] ), .ip2(n17641), .s(n17576), .op(n14302) );
  mux2_1 U20720 ( .ip1(\LUT[52][3] ), .ip2(n17642), .s(n17576), .op(n14301) );
  mux2_1 U20721 ( .ip1(\LUT[52][2] ), .ip2(n17643), .s(n17576), .op(n14300) );
  mux2_1 U20722 ( .ip1(\LUT[52][1] ), .ip2(n17644), .s(n17576), .op(n14299) );
  mux2_1 U20723 ( .ip1(\LUT[52][0] ), .ip2(n17646), .s(n17576), .op(n14298) );
  mux2_1 U20724 ( .ip1(\LUT[51][15] ), .ip2(d[15]), .s(n17577), .op(n14297) );
  mux2_1 U20725 ( .ip1(\LUT[51][14] ), .ip2(d[14]), .s(n17577), .op(n14296) );
  mux2_1 U20726 ( .ip1(\LUT[51][13] ), .ip2(d[13]), .s(n17577), .op(n14295) );
  mux2_1 U20727 ( .ip1(\LUT[51][12] ), .ip2(d[12]), .s(n17577), .op(n14294) );
  mux2_1 U20728 ( .ip1(\LUT[51][11] ), .ip2(d[11]), .s(n17577), .op(n14293) );
  mux2_1 U20729 ( .ip1(\LUT[51][10] ), .ip2(d[10]), .s(n17577), .op(n14292) );
  mux2_1 U20730 ( .ip1(\LUT[51][9] ), .ip2(d[9]), .s(n17577), .op(n14291) );
  mux2_1 U20731 ( .ip1(\LUT[51][8] ), .ip2(d[8]), .s(n17577), .op(n14290) );
  mux2_1 U20732 ( .ip1(\LUT[51][7] ), .ip2(d[7]), .s(n17577), .op(n14289) );
  mux2_1 U20733 ( .ip1(\LUT[51][6] ), .ip2(d[6]), .s(n17577), .op(n14288) );
  mux2_1 U20734 ( .ip1(\LUT[51][5] ), .ip2(d[5]), .s(n17578), .op(n14287) );
  mux2_1 U20735 ( .ip1(\LUT[51][4] ), .ip2(d[4]), .s(n17578), .op(n14286) );
  mux2_1 U20736 ( .ip1(\LUT[51][3] ), .ip2(d[3]), .s(n17578), .op(n14285) );
  mux2_1 U20737 ( .ip1(\LUT[51][2] ), .ip2(d[2]), .s(n17578), .op(n14284) );
  mux2_1 U20738 ( .ip1(\LUT[51][1] ), .ip2(d[1]), .s(n17578), .op(n14283) );
  mux2_1 U20739 ( .ip1(\LUT[51][0] ), .ip2(d[0]), .s(n17578), .op(n14282) );
  mux2_1 U20740 ( .ip1(\LUT[50][15] ), .ip2(n17629), .s(n17579), .op(n14281)
         );
  mux2_1 U20741 ( .ip1(\LUT[50][14] ), .ip2(n17630), .s(n17579), .op(n14280)
         );
  mux2_1 U20742 ( .ip1(\LUT[50][13] ), .ip2(n17631), .s(n17579), .op(n14279)
         );
  mux2_1 U20743 ( .ip1(\LUT[50][12] ), .ip2(n17632), .s(n17579), .op(n14278)
         );
  mux2_1 U20744 ( .ip1(\LUT[50][11] ), .ip2(n17633), .s(n17579), .op(n14277)
         );
  mux2_1 U20745 ( .ip1(\LUT[50][10] ), .ip2(n17634), .s(n17579), .op(n14276)
         );
  mux2_1 U20746 ( .ip1(\LUT[50][9] ), .ip2(n17635), .s(n17579), .op(n14275) );
  mux2_1 U20747 ( .ip1(\LUT[50][8] ), .ip2(n17636), .s(n17579), .op(n14274) );
  mux2_1 U20748 ( .ip1(\LUT[50][7] ), .ip2(n17637), .s(n17579), .op(n14273) );
  mux2_1 U20749 ( .ip1(\LUT[50][6] ), .ip2(n17639), .s(n17579), .op(n14272) );
  mux2_1 U20750 ( .ip1(\LUT[50][5] ), .ip2(n17640), .s(n17580), .op(n14271) );
  mux2_1 U20751 ( .ip1(\LUT[50][4] ), .ip2(n17641), .s(n17580), .op(n14270) );
  mux2_1 U20752 ( .ip1(\LUT[50][3] ), .ip2(n17642), .s(n17580), .op(n14269) );
  mux2_1 U20753 ( .ip1(\LUT[50][2] ), .ip2(n17643), .s(n17580), .op(n14268) );
  mux2_1 U20754 ( .ip1(\LUT[50][1] ), .ip2(n17644), .s(n17580), .op(n14267) );
  mux2_1 U20755 ( .ip1(\LUT[50][0] ), .ip2(n17646), .s(n17580), .op(n14266) );
  mux2_1 U20756 ( .ip1(\LUT[49][15] ), .ip2(d[15]), .s(n17581), .op(n14265) );
  mux2_1 U20757 ( .ip1(\LUT[49][14] ), .ip2(d[14]), .s(n17581), .op(n14264) );
  mux2_1 U20758 ( .ip1(\LUT[49][13] ), .ip2(d[13]), .s(n17581), .op(n14263) );
  mux2_1 U20759 ( .ip1(\LUT[49][12] ), .ip2(d[12]), .s(n17581), .op(n14262) );
  mux2_1 U20760 ( .ip1(\LUT[49][11] ), .ip2(d[11]), .s(n17581), .op(n14261) );
  mux2_1 U20761 ( .ip1(\LUT[49][10] ), .ip2(d[10]), .s(n17581), .op(n14260) );
  mux2_1 U20762 ( .ip1(\LUT[49][9] ), .ip2(d[9]), .s(n17581), .op(n14259) );
  mux2_1 U20763 ( .ip1(\LUT[49][8] ), .ip2(d[8]), .s(n17581), .op(n14258) );
  mux2_1 U20764 ( .ip1(\LUT[49][7] ), .ip2(d[7]), .s(n17581), .op(n14257) );
  mux2_1 U20765 ( .ip1(\LUT[49][6] ), .ip2(d[6]), .s(n17581), .op(n14256) );
  mux2_1 U20766 ( .ip1(\LUT[49][5] ), .ip2(d[5]), .s(n17582), .op(n14255) );
  mux2_1 U20767 ( .ip1(\LUT[49][4] ), .ip2(d[4]), .s(n17582), .op(n14254) );
  mux2_1 U20768 ( .ip1(\LUT[49][3] ), .ip2(d[3]), .s(n17582), .op(n14253) );
  mux2_1 U20769 ( .ip1(\LUT[49][2] ), .ip2(d[2]), .s(n17582), .op(n14252) );
  mux2_1 U20770 ( .ip1(\LUT[49][1] ), .ip2(d[1]), .s(n17582), .op(n14251) );
  mux2_1 U20771 ( .ip1(\LUT[49][0] ), .ip2(d[0]), .s(n17582), .op(n14250) );
  mux2_1 U20772 ( .ip1(\LUT[48][15] ), .ip2(n17629), .s(n17583), .op(n14249)
         );
  mux2_1 U20773 ( .ip1(\LUT[48][14] ), .ip2(n17630), .s(n17583), .op(n14248)
         );
  mux2_1 U20774 ( .ip1(\LUT[48][13] ), .ip2(n17631), .s(n17583), .op(n14247)
         );
  mux2_1 U20775 ( .ip1(\LUT[48][12] ), .ip2(n17632), .s(n17583), .op(n14246)
         );
  mux2_1 U20776 ( .ip1(\LUT[48][11] ), .ip2(n17633), .s(n17583), .op(n14245)
         );
  mux2_1 U20777 ( .ip1(\LUT[48][10] ), .ip2(n17634), .s(n17583), .op(n14244)
         );
  mux2_1 U20778 ( .ip1(\LUT[48][9] ), .ip2(n17635), .s(n17583), .op(n14243) );
  mux2_1 U20779 ( .ip1(\LUT[48][8] ), .ip2(n17636), .s(n17583), .op(n14242) );
  mux2_1 U20780 ( .ip1(\LUT[48][7] ), .ip2(n17637), .s(n17583), .op(n14241) );
  mux2_1 U20781 ( .ip1(\LUT[48][6] ), .ip2(n17639), .s(n17583), .op(n14240) );
  mux2_1 U20782 ( .ip1(\LUT[48][5] ), .ip2(n17640), .s(n17584), .op(n14239) );
  mux2_1 U20783 ( .ip1(\LUT[48][4] ), .ip2(n17641), .s(n17584), .op(n14238) );
  mux2_1 U20784 ( .ip1(\LUT[48][3] ), .ip2(n17642), .s(n17584), .op(n14237) );
  mux2_1 U20785 ( .ip1(\LUT[48][2] ), .ip2(n17643), .s(n17584), .op(n14236) );
  mux2_1 U20786 ( .ip1(\LUT[48][1] ), .ip2(n17644), .s(n17584), .op(n14235) );
  mux2_1 U20787 ( .ip1(\LUT[48][0] ), .ip2(n17646), .s(n17584), .op(n14234) );
  mux2_1 U20788 ( .ip1(\LUT[47][15] ), .ip2(n17629), .s(n17585), .op(n14233)
         );
  mux2_1 U20789 ( .ip1(\LUT[47][14] ), .ip2(n17630), .s(n17585), .op(n14232)
         );
  mux2_1 U20790 ( .ip1(\LUT[47][13] ), .ip2(n17631), .s(n17585), .op(n14231)
         );
  mux2_1 U20791 ( .ip1(\LUT[47][12] ), .ip2(n17632), .s(n17585), .op(n14230)
         );
  mux2_1 U20792 ( .ip1(\LUT[47][11] ), .ip2(n17633), .s(n17585), .op(n14229)
         );
  mux2_1 U20793 ( .ip1(\LUT[47][10] ), .ip2(n17634), .s(n17585), .op(n14228)
         );
  mux2_1 U20794 ( .ip1(\LUT[47][9] ), .ip2(n17635), .s(n17585), .op(n14227) );
  mux2_1 U20795 ( .ip1(\LUT[47][8] ), .ip2(n17636), .s(n17585), .op(n14226) );
  mux2_1 U20796 ( .ip1(\LUT[47][7] ), .ip2(n17637), .s(n17585), .op(n14225) );
  mux2_1 U20797 ( .ip1(\LUT[47][6] ), .ip2(n17639), .s(n17585), .op(n14224) );
  mux2_1 U20798 ( .ip1(\LUT[47][5] ), .ip2(n17640), .s(n17586), .op(n14223) );
  mux2_1 U20799 ( .ip1(\LUT[47][4] ), .ip2(n17641), .s(n17586), .op(n14222) );
  mux2_1 U20800 ( .ip1(\LUT[47][3] ), .ip2(n17642), .s(n17586), .op(n14221) );
  mux2_1 U20801 ( .ip1(\LUT[47][2] ), .ip2(n17643), .s(n17586), .op(n14220) );
  mux2_1 U20802 ( .ip1(\LUT[47][1] ), .ip2(n17644), .s(n17586), .op(n14219) );
  mux2_1 U20803 ( .ip1(\LUT[47][0] ), .ip2(n17646), .s(n17586), .op(n14218) );
  mux2_1 U20804 ( .ip1(\LUT[46][15] ), .ip2(n17629), .s(n17587), .op(n14217)
         );
  mux2_1 U20805 ( .ip1(\LUT[46][14] ), .ip2(n17630), .s(n17587), .op(n14216)
         );
  mux2_1 U20806 ( .ip1(\LUT[46][13] ), .ip2(n17631), .s(n17587), .op(n14215)
         );
  mux2_1 U20807 ( .ip1(\LUT[46][12] ), .ip2(n17632), .s(n17587), .op(n14214)
         );
  mux2_1 U20808 ( .ip1(\LUT[46][11] ), .ip2(n17633), .s(n17587), .op(n14213)
         );
  mux2_1 U20809 ( .ip1(\LUT[46][10] ), .ip2(n17634), .s(n17587), .op(n14212)
         );
  mux2_1 U20810 ( .ip1(\LUT[46][9] ), .ip2(n17635), .s(n17587), .op(n14211) );
  mux2_1 U20811 ( .ip1(\LUT[46][8] ), .ip2(n17636), .s(n17587), .op(n14210) );
  mux2_1 U20812 ( .ip1(\LUT[46][7] ), .ip2(n17637), .s(n17587), .op(n14209) );
  mux2_1 U20813 ( .ip1(\LUT[46][6] ), .ip2(n17639), .s(n17587), .op(n14208) );
  mux2_1 U20814 ( .ip1(\LUT[46][5] ), .ip2(n17640), .s(n17588), .op(n14207) );
  mux2_1 U20815 ( .ip1(\LUT[46][4] ), .ip2(n17641), .s(n17588), .op(n14206) );
  mux2_1 U20816 ( .ip1(\LUT[46][3] ), .ip2(n17642), .s(n17588), .op(n14205) );
  mux2_1 U20817 ( .ip1(\LUT[46][2] ), .ip2(n17643), .s(n17588), .op(n14204) );
  mux2_1 U20818 ( .ip1(\LUT[46][1] ), .ip2(n17644), .s(n17588), .op(n14203) );
  mux2_1 U20819 ( .ip1(\LUT[46][0] ), .ip2(n17646), .s(n17588), .op(n14202) );
  mux2_1 U20820 ( .ip1(\LUT[45][15] ), .ip2(n17629), .s(n17589), .op(n14201)
         );
  mux2_1 U20821 ( .ip1(\LUT[45][14] ), .ip2(n17630), .s(n17589), .op(n14200)
         );
  mux2_1 U20822 ( .ip1(\LUT[45][13] ), .ip2(n17631), .s(n17589), .op(n14199)
         );
  mux2_1 U20823 ( .ip1(\LUT[45][12] ), .ip2(n17632), .s(n17589), .op(n14198)
         );
  mux2_1 U20824 ( .ip1(\LUT[45][11] ), .ip2(n17633), .s(n17589), .op(n14197)
         );
  mux2_1 U20825 ( .ip1(\LUT[45][10] ), .ip2(n17634), .s(n17589), .op(n14196)
         );
  mux2_1 U20826 ( .ip1(\LUT[45][9] ), .ip2(n17635), .s(n17589), .op(n14195) );
  mux2_1 U20827 ( .ip1(\LUT[45][8] ), .ip2(n17636), .s(n17589), .op(n14194) );
  mux2_1 U20828 ( .ip1(\LUT[45][7] ), .ip2(n17637), .s(n17589), .op(n14193) );
  mux2_1 U20829 ( .ip1(\LUT[45][6] ), .ip2(n17639), .s(n17589), .op(n14192) );
  mux2_1 U20830 ( .ip1(\LUT[45][5] ), .ip2(n17640), .s(n17590), .op(n14191) );
  mux2_1 U20831 ( .ip1(\LUT[45][4] ), .ip2(n17641), .s(n17590), .op(n14190) );
  mux2_1 U20832 ( .ip1(\LUT[45][3] ), .ip2(n17642), .s(n17590), .op(n14189) );
  mux2_1 U20833 ( .ip1(\LUT[45][2] ), .ip2(n17643), .s(n17590), .op(n14188) );
  mux2_1 U20834 ( .ip1(\LUT[45][1] ), .ip2(n17644), .s(n17590), .op(n14187) );
  mux2_1 U20835 ( .ip1(\LUT[45][0] ), .ip2(n17646), .s(n17590), .op(n14186) );
  mux2_1 U20836 ( .ip1(\LUT[44][15] ), .ip2(n17629), .s(n17591), .op(n14185)
         );
  mux2_1 U20837 ( .ip1(\LUT[44][14] ), .ip2(n17630), .s(n17591), .op(n14184)
         );
  mux2_1 U20838 ( .ip1(\LUT[44][13] ), .ip2(n17631), .s(n17591), .op(n14183)
         );
  mux2_1 U20839 ( .ip1(\LUT[44][12] ), .ip2(n17632), .s(n17591), .op(n14182)
         );
  mux2_1 U20840 ( .ip1(\LUT[44][11] ), .ip2(n17633), .s(n17591), .op(n14181)
         );
  mux2_1 U20841 ( .ip1(\LUT[44][10] ), .ip2(n17634), .s(n17591), .op(n14180)
         );
  mux2_1 U20842 ( .ip1(\LUT[44][9] ), .ip2(n17635), .s(n17591), .op(n14179) );
  mux2_1 U20843 ( .ip1(\LUT[44][8] ), .ip2(n17636), .s(n17591), .op(n14178) );
  mux2_1 U20844 ( .ip1(\LUT[44][7] ), .ip2(n17637), .s(n17591), .op(n14177) );
  mux2_1 U20845 ( .ip1(\LUT[44][6] ), .ip2(n17639), .s(n17591), .op(n14176) );
  mux2_1 U20846 ( .ip1(\LUT[44][5] ), .ip2(n17640), .s(n17592), .op(n14175) );
  mux2_1 U20847 ( .ip1(\LUT[44][4] ), .ip2(n17641), .s(n17592), .op(n14174) );
  mux2_1 U20848 ( .ip1(\LUT[44][3] ), .ip2(n17642), .s(n17592), .op(n14173) );
  mux2_1 U20849 ( .ip1(\LUT[44][2] ), .ip2(n17643), .s(n17592), .op(n14172) );
  mux2_1 U20850 ( .ip1(\LUT[44][1] ), .ip2(n17644), .s(n17592), .op(n14171) );
  mux2_1 U20851 ( .ip1(\LUT[44][0] ), .ip2(n17646), .s(n17592), .op(n14170) );
  mux2_1 U20852 ( .ip1(\LUT[43][15] ), .ip2(n17629), .s(n17593), .op(n14169)
         );
  mux2_1 U20853 ( .ip1(\LUT[43][14] ), .ip2(n17630), .s(n17593), .op(n14168)
         );
  mux2_1 U20854 ( .ip1(\LUT[43][13] ), .ip2(n17631), .s(n17593), .op(n14167)
         );
  mux2_1 U20855 ( .ip1(\LUT[43][12] ), .ip2(n17632), .s(n17593), .op(n14166)
         );
  mux2_1 U20856 ( .ip1(\LUT[43][11] ), .ip2(n17633), .s(n17593), .op(n14165)
         );
  mux2_1 U20857 ( .ip1(\LUT[43][10] ), .ip2(n17634), .s(n17593), .op(n14164)
         );
  mux2_1 U20858 ( .ip1(\LUT[43][9] ), .ip2(n17635), .s(n17593), .op(n14163) );
  mux2_1 U20859 ( .ip1(\LUT[43][8] ), .ip2(n17636), .s(n17593), .op(n14162) );
  mux2_1 U20860 ( .ip1(\LUT[43][7] ), .ip2(n17637), .s(n17593), .op(n14161) );
  mux2_1 U20861 ( .ip1(\LUT[43][6] ), .ip2(n17639), .s(n17593), .op(n14160) );
  mux2_1 U20862 ( .ip1(\LUT[43][5] ), .ip2(n17640), .s(n17594), .op(n14159) );
  mux2_1 U20863 ( .ip1(\LUT[43][4] ), .ip2(n17641), .s(n17594), .op(n14158) );
  mux2_1 U20864 ( .ip1(\LUT[43][3] ), .ip2(n17642), .s(n17594), .op(n14157) );
  mux2_1 U20865 ( .ip1(\LUT[43][2] ), .ip2(n17643), .s(n17594), .op(n14156) );
  mux2_1 U20866 ( .ip1(\LUT[43][1] ), .ip2(n17644), .s(n17594), .op(n14155) );
  mux2_1 U20867 ( .ip1(\LUT[43][0] ), .ip2(n17646), .s(n17594), .op(n14154) );
  mux2_1 U20868 ( .ip1(\LUT[42][15] ), .ip2(d[15]), .s(n17595), .op(n14153) );
  mux2_1 U20869 ( .ip1(\LUT[42][14] ), .ip2(d[14]), .s(n17595), .op(n14152) );
  mux2_1 U20870 ( .ip1(\LUT[42][13] ), .ip2(d[13]), .s(n17595), .op(n14151) );
  mux2_1 U20871 ( .ip1(\LUT[42][12] ), .ip2(d[12]), .s(n17595), .op(n14150) );
  mux2_1 U20872 ( .ip1(\LUT[42][11] ), .ip2(d[11]), .s(n17595), .op(n14149) );
  mux2_1 U20873 ( .ip1(\LUT[42][10] ), .ip2(d[10]), .s(n17595), .op(n14148) );
  mux2_1 U20874 ( .ip1(\LUT[42][9] ), .ip2(d[9]), .s(n17595), .op(n14147) );
  mux2_1 U20875 ( .ip1(\LUT[42][8] ), .ip2(d[8]), .s(n17595), .op(n14146) );
  mux2_1 U20876 ( .ip1(\LUT[42][7] ), .ip2(d[7]), .s(n17595), .op(n14145) );
  mux2_1 U20877 ( .ip1(\LUT[42][6] ), .ip2(d[6]), .s(n17595), .op(n14144) );
  mux2_1 U20878 ( .ip1(\LUT[42][5] ), .ip2(d[5]), .s(n17596), .op(n14143) );
  mux2_1 U20879 ( .ip1(\LUT[42][4] ), .ip2(d[4]), .s(n17596), .op(n14142) );
  mux2_1 U20880 ( .ip1(\LUT[42][3] ), .ip2(d[3]), .s(n17596), .op(n14141) );
  mux2_1 U20881 ( .ip1(\LUT[42][2] ), .ip2(d[2]), .s(n17596), .op(n14140) );
  mux2_1 U20882 ( .ip1(\LUT[42][1] ), .ip2(d[1]), .s(n17596), .op(n14139) );
  mux2_1 U20883 ( .ip1(\LUT[42][0] ), .ip2(d[0]), .s(n17596), .op(n14138) );
  mux2_1 U20884 ( .ip1(\LUT[41][15] ), .ip2(n17629), .s(n17597), .op(n14137)
         );
  mux2_1 U20885 ( .ip1(\LUT[41][14] ), .ip2(n17630), .s(n17597), .op(n14136)
         );
  mux2_1 U20886 ( .ip1(\LUT[41][13] ), .ip2(n17631), .s(n17597), .op(n14135)
         );
  mux2_1 U20887 ( .ip1(\LUT[41][12] ), .ip2(n17632), .s(n17597), .op(n14134)
         );
  mux2_1 U20888 ( .ip1(\LUT[41][11] ), .ip2(n17633), .s(n17597), .op(n14133)
         );
  mux2_1 U20889 ( .ip1(\LUT[41][10] ), .ip2(n17634), .s(n17597), .op(n14132)
         );
  mux2_1 U20890 ( .ip1(\LUT[41][9] ), .ip2(n17635), .s(n17597), .op(n14131) );
  mux2_1 U20891 ( .ip1(\LUT[41][8] ), .ip2(n17636), .s(n17597), .op(n14130) );
  mux2_1 U20892 ( .ip1(\LUT[41][7] ), .ip2(n17637), .s(n17597), .op(n14129) );
  mux2_1 U20893 ( .ip1(\LUT[41][6] ), .ip2(n17639), .s(n17597), .op(n14128) );
  mux2_1 U20894 ( .ip1(\LUT[41][5] ), .ip2(n17640), .s(n17598), .op(n14127) );
  mux2_1 U20895 ( .ip1(\LUT[41][4] ), .ip2(n17641), .s(n17598), .op(n14126) );
  mux2_1 U20896 ( .ip1(\LUT[41][3] ), .ip2(n17642), .s(n17598), .op(n14125) );
  mux2_1 U20897 ( .ip1(\LUT[41][2] ), .ip2(n17643), .s(n17598), .op(n14124) );
  mux2_1 U20898 ( .ip1(\LUT[41][1] ), .ip2(n17644), .s(n17598), .op(n14123) );
  mux2_1 U20899 ( .ip1(\LUT[41][0] ), .ip2(n17646), .s(n17598), .op(n14122) );
  mux2_1 U20900 ( .ip1(\LUT[40][15] ), .ip2(d[15]), .s(n17599), .op(n14121) );
  mux2_1 U20901 ( .ip1(\LUT[40][14] ), .ip2(d[14]), .s(n17599), .op(n14120) );
  mux2_1 U20902 ( .ip1(\LUT[40][13] ), .ip2(d[13]), .s(n17599), .op(n14119) );
  mux2_1 U20903 ( .ip1(\LUT[40][12] ), .ip2(d[12]), .s(n17599), .op(n14118) );
  mux2_1 U20904 ( .ip1(\LUT[40][11] ), .ip2(d[11]), .s(n17599), .op(n14117) );
  mux2_1 U20905 ( .ip1(\LUT[40][10] ), .ip2(d[10]), .s(n17599), .op(n14116) );
  mux2_1 U20906 ( .ip1(\LUT[40][9] ), .ip2(d[9]), .s(n17599), .op(n14115) );
  mux2_1 U20907 ( .ip1(\LUT[40][8] ), .ip2(d[8]), .s(n17599), .op(n14114) );
  mux2_1 U20908 ( .ip1(\LUT[40][7] ), .ip2(d[7]), .s(n17599), .op(n14113) );
  mux2_1 U20909 ( .ip1(\LUT[40][6] ), .ip2(d[6]), .s(n17599), .op(n14112) );
  mux2_1 U20910 ( .ip1(\LUT[40][5] ), .ip2(d[5]), .s(n17600), .op(n14111) );
  mux2_1 U20911 ( .ip1(\LUT[40][4] ), .ip2(d[4]), .s(n17600), .op(n14110) );
  mux2_1 U20912 ( .ip1(\LUT[40][3] ), .ip2(d[3]), .s(n17600), .op(n14109) );
  mux2_1 U20913 ( .ip1(\LUT[40][2] ), .ip2(d[2]), .s(n17600), .op(n14108) );
  mux2_1 U20914 ( .ip1(\LUT[40][1] ), .ip2(d[1]), .s(n17600), .op(n14107) );
  mux2_1 U20915 ( .ip1(\LUT[40][0] ), .ip2(d[0]), .s(n17600), .op(n14106) );
  mux2_1 U20916 ( .ip1(\LUT[39][15] ), .ip2(n17629), .s(n17601), .op(n14105)
         );
  mux2_1 U20917 ( .ip1(\LUT[39][14] ), .ip2(n17630), .s(n17601), .op(n14104)
         );
  mux2_1 U20918 ( .ip1(\LUT[39][13] ), .ip2(n17631), .s(n17601), .op(n14103)
         );
  mux2_1 U20919 ( .ip1(\LUT[39][12] ), .ip2(n17632), .s(n17601), .op(n14102)
         );
  mux2_1 U20920 ( .ip1(\LUT[39][11] ), .ip2(n17633), .s(n17601), .op(n14101)
         );
  mux2_1 U20921 ( .ip1(\LUT[39][10] ), .ip2(n17634), .s(n17601), .op(n14100)
         );
  mux2_1 U20922 ( .ip1(\LUT[39][9] ), .ip2(n17635), .s(n17601), .op(n14099) );
  mux2_1 U20923 ( .ip1(\LUT[39][8] ), .ip2(n17636), .s(n17601), .op(n14098) );
  mux2_1 U20924 ( .ip1(\LUT[39][7] ), .ip2(n17637), .s(n17601), .op(n14097) );
  mux2_1 U20925 ( .ip1(\LUT[39][6] ), .ip2(n17639), .s(n17601), .op(n14096) );
  mux2_1 U20926 ( .ip1(\LUT[39][5] ), .ip2(n17640), .s(n17602), .op(n14095) );
  mux2_1 U20927 ( .ip1(\LUT[39][4] ), .ip2(n17641), .s(n17602), .op(n14094) );
  mux2_1 U20928 ( .ip1(\LUT[39][3] ), .ip2(n17642), .s(n17602), .op(n14093) );
  mux2_1 U20929 ( .ip1(\LUT[39][2] ), .ip2(n17643), .s(n17602), .op(n14092) );
  mux2_1 U20930 ( .ip1(\LUT[39][1] ), .ip2(n17644), .s(n17602), .op(n14091) );
  mux2_1 U20931 ( .ip1(\LUT[39][0] ), .ip2(n17646), .s(n17602), .op(n14090) );
  mux2_1 U20932 ( .ip1(\LUT[38][15] ), .ip2(n17629), .s(n17603), .op(n14089)
         );
  mux2_1 U20933 ( .ip1(\LUT[38][14] ), .ip2(n17630), .s(n17603), .op(n14088)
         );
  mux2_1 U20934 ( .ip1(\LUT[38][13] ), .ip2(n17631), .s(n17603), .op(n14087)
         );
  mux2_1 U20935 ( .ip1(\LUT[38][12] ), .ip2(n17632), .s(n17603), .op(n14086)
         );
  mux2_1 U20936 ( .ip1(\LUT[38][11] ), .ip2(n17633), .s(n17603), .op(n14085)
         );
  mux2_1 U20937 ( .ip1(\LUT[38][10] ), .ip2(n17634), .s(n17603), .op(n14084)
         );
  mux2_1 U20938 ( .ip1(\LUT[38][9] ), .ip2(n17635), .s(n17603), .op(n14083) );
  mux2_1 U20939 ( .ip1(\LUT[38][8] ), .ip2(n17636), .s(n17603), .op(n14082) );
  mux2_1 U20940 ( .ip1(\LUT[38][7] ), .ip2(n17637), .s(n17603), .op(n14081) );
  mux2_1 U20941 ( .ip1(\LUT[38][6] ), .ip2(n17639), .s(n17603), .op(n14080) );
  mux2_1 U20942 ( .ip1(\LUT[38][5] ), .ip2(n17640), .s(n17604), .op(n14079) );
  mux2_1 U20943 ( .ip1(\LUT[38][4] ), .ip2(n17641), .s(n17604), .op(n14078) );
  mux2_1 U20944 ( .ip1(\LUT[38][3] ), .ip2(n17642), .s(n17604), .op(n14077) );
  mux2_1 U20945 ( .ip1(\LUT[38][2] ), .ip2(n17643), .s(n17604), .op(n14076) );
  mux2_1 U20946 ( .ip1(\LUT[38][1] ), .ip2(n17644), .s(n17604), .op(n14075) );
  mux2_1 U20947 ( .ip1(\LUT[38][0] ), .ip2(n17646), .s(n17604), .op(n14074) );
  mux2_1 U20948 ( .ip1(\LUT[37][15] ), .ip2(n17629), .s(n17605), .op(n14073)
         );
  mux2_1 U20949 ( .ip1(\LUT[37][14] ), .ip2(n17630), .s(n17605), .op(n14072)
         );
  mux2_1 U20950 ( .ip1(\LUT[37][13] ), .ip2(n17631), .s(n17605), .op(n14071)
         );
  mux2_1 U20951 ( .ip1(\LUT[37][12] ), .ip2(n17632), .s(n17605), .op(n14070)
         );
  mux2_1 U20952 ( .ip1(\LUT[37][11] ), .ip2(n17633), .s(n17605), .op(n14069)
         );
  mux2_1 U20953 ( .ip1(\LUT[37][10] ), .ip2(n17634), .s(n17605), .op(n14068)
         );
  mux2_1 U20954 ( .ip1(\LUT[37][9] ), .ip2(n17635), .s(n17605), .op(n14067) );
  mux2_1 U20955 ( .ip1(\LUT[37][8] ), .ip2(n17636), .s(n17605), .op(n14066) );
  mux2_1 U20956 ( .ip1(\LUT[37][7] ), .ip2(n17637), .s(n17605), .op(n14065) );
  mux2_1 U20957 ( .ip1(\LUT[37][6] ), .ip2(n17639), .s(n17605), .op(n14064) );
  mux2_1 U20958 ( .ip1(\LUT[37][5] ), .ip2(n17640), .s(n17606), .op(n14063) );
  mux2_1 U20959 ( .ip1(\LUT[37][4] ), .ip2(n17641), .s(n17606), .op(n14062) );
  mux2_1 U20960 ( .ip1(\LUT[37][3] ), .ip2(n17642), .s(n17606), .op(n14061) );
  mux2_1 U20961 ( .ip1(\LUT[37][2] ), .ip2(n17643), .s(n17606), .op(n14060) );
  mux2_1 U20962 ( .ip1(\LUT[37][1] ), .ip2(n17644), .s(n17606), .op(n14059) );
  mux2_1 U20963 ( .ip1(\LUT[37][0] ), .ip2(n17646), .s(n17606), .op(n14058) );
  mux2_1 U20964 ( .ip1(\LUT[36][15] ), .ip2(d[15]), .s(n17607), .op(n14057) );
  mux2_1 U20965 ( .ip1(\LUT[36][14] ), .ip2(d[14]), .s(n17607), .op(n14056) );
  mux2_1 U20966 ( .ip1(\LUT[36][13] ), .ip2(d[13]), .s(n17607), .op(n14055) );
  mux2_1 U20967 ( .ip1(\LUT[36][12] ), .ip2(d[12]), .s(n17607), .op(n14054) );
  mux2_1 U20968 ( .ip1(\LUT[36][11] ), .ip2(d[11]), .s(n17607), .op(n14053) );
  mux2_1 U20969 ( .ip1(\LUT[36][10] ), .ip2(d[10]), .s(n17607), .op(n14052) );
  mux2_1 U20970 ( .ip1(\LUT[36][9] ), .ip2(d[9]), .s(n17607), .op(n14051) );
  mux2_1 U20971 ( .ip1(\LUT[36][8] ), .ip2(d[8]), .s(n17607), .op(n14050) );
  mux2_1 U20972 ( .ip1(\LUT[36][7] ), .ip2(d[7]), .s(n17607), .op(n14049) );
  mux2_1 U20973 ( .ip1(\LUT[36][6] ), .ip2(d[6]), .s(n17607), .op(n14048) );
  mux2_1 U20974 ( .ip1(\LUT[36][5] ), .ip2(d[5]), .s(n17608), .op(n14047) );
  mux2_1 U20975 ( .ip1(\LUT[36][4] ), .ip2(d[4]), .s(n17608), .op(n14046) );
  mux2_1 U20976 ( .ip1(\LUT[36][3] ), .ip2(d[3]), .s(n17608), .op(n14045) );
  mux2_1 U20977 ( .ip1(\LUT[36][2] ), .ip2(d[2]), .s(n17608), .op(n14044) );
  mux2_1 U20978 ( .ip1(\LUT[36][1] ), .ip2(d[1]), .s(n17608), .op(n14043) );
  mux2_1 U20979 ( .ip1(\LUT[36][0] ), .ip2(d[0]), .s(n17608), .op(n14042) );
  mux2_1 U20980 ( .ip1(\LUT[35][15] ), .ip2(n17629), .s(n17609), .op(n14041)
         );
  mux2_1 U20981 ( .ip1(\LUT[35][14] ), .ip2(n17630), .s(n17609), .op(n14040)
         );
  mux2_1 U20982 ( .ip1(\LUT[35][13] ), .ip2(n17631), .s(n17609), .op(n14039)
         );
  mux2_1 U20983 ( .ip1(\LUT[35][12] ), .ip2(n17632), .s(n17609), .op(n14038)
         );
  mux2_1 U20984 ( .ip1(\LUT[35][11] ), .ip2(n17633), .s(n17609), .op(n14037)
         );
  mux2_1 U20985 ( .ip1(\LUT[35][10] ), .ip2(n17634), .s(n17609), .op(n14036)
         );
  mux2_1 U20986 ( .ip1(\LUT[35][9] ), .ip2(n17635), .s(n17609), .op(n14035) );
  mux2_1 U20987 ( .ip1(\LUT[35][8] ), .ip2(n17636), .s(n17609), .op(n14034) );
  mux2_1 U20988 ( .ip1(\LUT[35][7] ), .ip2(n17637), .s(n17609), .op(n14033) );
  mux2_1 U20989 ( .ip1(\LUT[35][6] ), .ip2(n17639), .s(n17609), .op(n14032) );
  mux2_1 U20990 ( .ip1(\LUT[35][5] ), .ip2(n17640), .s(n17610), .op(n14031) );
  mux2_1 U20991 ( .ip1(\LUT[35][4] ), .ip2(n17641), .s(n17610), .op(n14030) );
  mux2_1 U20992 ( .ip1(\LUT[35][3] ), .ip2(n17642), .s(n17610), .op(n14029) );
  mux2_1 U20993 ( .ip1(\LUT[35][2] ), .ip2(n17643), .s(n17610), .op(n14028) );
  mux2_1 U20994 ( .ip1(\LUT[35][1] ), .ip2(n17644), .s(n17610), .op(n14027) );
  mux2_1 U20995 ( .ip1(\LUT[35][0] ), .ip2(n17646), .s(n17610), .op(n14026) );
  mux2_1 U20996 ( .ip1(\LUT[34][15] ), .ip2(d[15]), .s(n17611), .op(n14025) );
  mux2_1 U20997 ( .ip1(\LUT[34][14] ), .ip2(d[14]), .s(n17611), .op(n14024) );
  mux2_1 U20998 ( .ip1(\LUT[34][13] ), .ip2(d[13]), .s(n17611), .op(n14023) );
  mux2_1 U20999 ( .ip1(\LUT[34][12] ), .ip2(d[12]), .s(n17611), .op(n14022) );
  mux2_1 U21000 ( .ip1(\LUT[34][11] ), .ip2(d[11]), .s(n17611), .op(n14021) );
  mux2_1 U21001 ( .ip1(\LUT[34][10] ), .ip2(d[10]), .s(n17611), .op(n14020) );
  mux2_1 U21002 ( .ip1(\LUT[34][9] ), .ip2(d[9]), .s(n17611), .op(n14019) );
  mux2_1 U21003 ( .ip1(\LUT[34][8] ), .ip2(d[8]), .s(n17611), .op(n14018) );
  mux2_1 U21004 ( .ip1(\LUT[34][7] ), .ip2(d[7]), .s(n17611), .op(n14017) );
  mux2_1 U21005 ( .ip1(\LUT[34][6] ), .ip2(d[6]), .s(n17611), .op(n14016) );
  mux2_1 U21006 ( .ip1(\LUT[34][5] ), .ip2(d[5]), .s(n17612), .op(n14015) );
  mux2_1 U21007 ( .ip1(\LUT[34][4] ), .ip2(d[4]), .s(n17612), .op(n14014) );
  mux2_1 U21008 ( .ip1(\LUT[34][3] ), .ip2(d[3]), .s(n17612), .op(n14013) );
  mux2_1 U21009 ( .ip1(\LUT[34][2] ), .ip2(d[2]), .s(n17612), .op(n14012) );
  mux2_1 U21010 ( .ip1(\LUT[34][1] ), .ip2(d[1]), .s(n17612), .op(n14011) );
  mux2_1 U21011 ( .ip1(\LUT[34][0] ), .ip2(d[0]), .s(n17612), .op(n14010) );
  mux2_1 U21012 ( .ip1(\LUT[33][15] ), .ip2(n17629), .s(n17613), .op(n14009)
         );
  mux2_1 U21013 ( .ip1(\LUT[33][14] ), .ip2(n17630), .s(n17613), .op(n14008)
         );
  mux2_1 U21014 ( .ip1(\LUT[33][13] ), .ip2(n17631), .s(n17613), .op(n14007)
         );
  mux2_1 U21015 ( .ip1(\LUT[33][12] ), .ip2(n17632), .s(n17613), .op(n14006)
         );
  mux2_1 U21016 ( .ip1(\LUT[33][11] ), .ip2(n17633), .s(n17613), .op(n14005)
         );
  mux2_1 U21017 ( .ip1(\LUT[33][10] ), .ip2(n17634), .s(n17613), .op(n14004)
         );
  mux2_1 U21018 ( .ip1(\LUT[33][9] ), .ip2(n17635), .s(n17613), .op(n14003) );
  mux2_1 U21019 ( .ip1(\LUT[33][8] ), .ip2(n17636), .s(n17613), .op(n14002) );
  mux2_1 U21020 ( .ip1(\LUT[33][7] ), .ip2(n17637), .s(n17613), .op(n14001) );
  mux2_1 U21021 ( .ip1(\LUT[33][6] ), .ip2(n17639), .s(n17613), .op(n14000) );
  mux2_1 U21022 ( .ip1(\LUT[33][5] ), .ip2(n17640), .s(n17614), .op(n13999) );
  mux2_1 U21023 ( .ip1(\LUT[33][4] ), .ip2(n17641), .s(n17614), .op(n13998) );
  mux2_1 U21024 ( .ip1(\LUT[33][3] ), .ip2(n17642), .s(n17614), .op(n13997) );
  mux2_1 U21025 ( .ip1(\LUT[33][2] ), .ip2(n17643), .s(n17614), .op(n13996) );
  mux2_1 U21026 ( .ip1(\LUT[33][1] ), .ip2(n17644), .s(n17614), .op(n13995) );
  mux2_1 U21027 ( .ip1(\LUT[33][0] ), .ip2(n17646), .s(n17614), .op(n13994) );
  mux2_1 U21028 ( .ip1(\LUT[32][15] ), .ip2(d[15]), .s(n17615), .op(n13993) );
  mux2_1 U21029 ( .ip1(\LUT[32][14] ), .ip2(d[14]), .s(n17615), .op(n13992) );
  mux2_1 U21030 ( .ip1(\LUT[32][13] ), .ip2(d[13]), .s(n17615), .op(n13991) );
  mux2_1 U21031 ( .ip1(\LUT[32][12] ), .ip2(d[12]), .s(n17615), .op(n13990) );
  mux2_1 U21032 ( .ip1(\LUT[32][11] ), .ip2(d[11]), .s(n17615), .op(n13989) );
  mux2_1 U21033 ( .ip1(\LUT[32][10] ), .ip2(d[10]), .s(n17615), .op(n13988) );
  mux2_1 U21034 ( .ip1(\LUT[32][9] ), .ip2(d[9]), .s(n17615), .op(n13987) );
  mux2_1 U21035 ( .ip1(\LUT[32][8] ), .ip2(d[8]), .s(n17615), .op(n13986) );
  mux2_1 U21036 ( .ip1(\LUT[32][7] ), .ip2(d[7]), .s(n17615), .op(n13985) );
  mux2_1 U21037 ( .ip1(\LUT[32][6] ), .ip2(d[6]), .s(n17615), .op(n13984) );
  mux2_1 U21038 ( .ip1(\LUT[32][5] ), .ip2(d[5]), .s(n17616), .op(n13983) );
  mux2_1 U21039 ( .ip1(\LUT[32][4] ), .ip2(d[4]), .s(n17616), .op(n13982) );
  mux2_1 U21040 ( .ip1(\LUT[32][3] ), .ip2(d[3]), .s(n17616), .op(n13981) );
  mux2_1 U21041 ( .ip1(\LUT[32][2] ), .ip2(d[2]), .s(n17616), .op(n13980) );
  mux2_1 U21042 ( .ip1(\LUT[32][1] ), .ip2(d[1]), .s(n17616), .op(n13979) );
  mux2_1 U21043 ( .ip1(\LUT[32][0] ), .ip2(d[0]), .s(n17616), .op(n13978) );
  mux2_1 U21044 ( .ip1(\LUT[31][15] ), .ip2(n17629), .s(n17617), .op(n13977)
         );
  mux2_1 U21045 ( .ip1(\LUT[31][14] ), .ip2(n17630), .s(n17617), .op(n13976)
         );
  mux2_1 U21046 ( .ip1(\LUT[31][13] ), .ip2(n17631), .s(n17617), .op(n13975)
         );
  mux2_1 U21047 ( .ip1(\LUT[31][12] ), .ip2(n17632), .s(n17617), .op(n13974)
         );
  mux2_1 U21048 ( .ip1(\LUT[31][11] ), .ip2(n17633), .s(n17617), .op(n13973)
         );
  mux2_1 U21049 ( .ip1(\LUT[31][10] ), .ip2(n17634), .s(n17617), .op(n13972)
         );
  mux2_1 U21050 ( .ip1(\LUT[31][9] ), .ip2(n17635), .s(n17617), .op(n13971) );
  mux2_1 U21051 ( .ip1(\LUT[31][8] ), .ip2(n17636), .s(n17617), .op(n13970) );
  mux2_1 U21052 ( .ip1(\LUT[31][7] ), .ip2(n17637), .s(n17617), .op(n13969) );
  mux2_1 U21053 ( .ip1(\LUT[31][6] ), .ip2(n17639), .s(n17617), .op(n13968) );
  mux2_1 U21054 ( .ip1(\LUT[31][5] ), .ip2(n17640), .s(n17618), .op(n13967) );
  mux2_1 U21055 ( .ip1(\LUT[31][4] ), .ip2(n17641), .s(n17618), .op(n13966) );
  mux2_1 U21056 ( .ip1(\LUT[31][3] ), .ip2(n17642), .s(n17618), .op(n13965) );
  mux2_1 U21057 ( .ip1(\LUT[31][2] ), .ip2(n17643), .s(n17618), .op(n13964) );
  mux2_1 U21058 ( .ip1(\LUT[31][1] ), .ip2(n17644), .s(n17618), .op(n13963) );
  mux2_1 U21059 ( .ip1(\LUT[31][0] ), .ip2(n17646), .s(n17618), .op(n13962) );
  mux2_1 U21060 ( .ip1(\LUT[30][15] ), .ip2(d[15]), .s(n17619), .op(n13961) );
  mux2_1 U21061 ( .ip1(\LUT[30][14] ), .ip2(d[14]), .s(n17619), .op(n13960) );
  mux2_1 U21062 ( .ip1(\LUT[30][13] ), .ip2(d[13]), .s(n17619), .op(n13959) );
  mux2_1 U21063 ( .ip1(\LUT[30][12] ), .ip2(d[12]), .s(n17619), .op(n13958) );
  mux2_1 U21064 ( .ip1(\LUT[30][11] ), .ip2(d[11]), .s(n17619), .op(n13957) );
  mux2_1 U21065 ( .ip1(\LUT[30][10] ), .ip2(d[10]), .s(n17619), .op(n13956) );
  mux2_1 U21066 ( .ip1(\LUT[30][9] ), .ip2(d[9]), .s(n17619), .op(n13955) );
  mux2_1 U21067 ( .ip1(\LUT[30][8] ), .ip2(d[8]), .s(n17619), .op(n13954) );
  mux2_1 U21068 ( .ip1(\LUT[30][7] ), .ip2(d[7]), .s(n17619), .op(n13953) );
  mux2_1 U21069 ( .ip1(\LUT[30][6] ), .ip2(d[6]), .s(n17619), .op(n13952) );
  mux2_1 U21070 ( .ip1(\LUT[30][5] ), .ip2(d[5]), .s(n17620), .op(n13951) );
  mux2_1 U21071 ( .ip1(\LUT[30][4] ), .ip2(d[4]), .s(n17620), .op(n13950) );
  mux2_1 U21072 ( .ip1(\LUT[30][3] ), .ip2(d[3]), .s(n17620), .op(n13949) );
  mux2_1 U21073 ( .ip1(\LUT[30][2] ), .ip2(d[2]), .s(n17620), .op(n13948) );
  mux2_1 U21074 ( .ip1(\LUT[30][1] ), .ip2(d[1]), .s(n17620), .op(n13947) );
  mux2_1 U21075 ( .ip1(\LUT[30][0] ), .ip2(d[0]), .s(n17620), .op(n13946) );
  mux2_1 U21076 ( .ip1(\LUT[29][15] ), .ip2(n17629), .s(n17621), .op(n13945)
         );
  mux2_1 U21077 ( .ip1(\LUT[29][14] ), .ip2(n17630), .s(n17621), .op(n13944)
         );
  mux2_1 U21078 ( .ip1(\LUT[29][13] ), .ip2(n17631), .s(n17621), .op(n13943)
         );
  mux2_1 U21079 ( .ip1(\LUT[29][12] ), .ip2(n17632), .s(n17621), .op(n13942)
         );
  mux2_1 U21080 ( .ip1(\LUT[29][11] ), .ip2(n17633), .s(n17621), .op(n13941)
         );
  mux2_1 U21081 ( .ip1(\LUT[29][10] ), .ip2(n17634), .s(n17621), .op(n13940)
         );
  mux2_1 U21082 ( .ip1(\LUT[29][9] ), .ip2(n17635), .s(n17621), .op(n13939) );
  mux2_1 U21083 ( .ip1(\LUT[29][8] ), .ip2(n17636), .s(n17621), .op(n13938) );
  mux2_1 U21084 ( .ip1(\LUT[29][7] ), .ip2(n17637), .s(n17621), .op(n13937) );
  mux2_1 U21085 ( .ip1(\LUT[29][6] ), .ip2(n17639), .s(n17621), .op(n13936) );
  mux2_1 U21086 ( .ip1(\LUT[29][5] ), .ip2(n17640), .s(n17622), .op(n13935) );
  mux2_1 U21087 ( .ip1(\LUT[29][4] ), .ip2(n17641), .s(n17622), .op(n13934) );
  mux2_1 U21088 ( .ip1(\LUT[29][3] ), .ip2(n17642), .s(n17622), .op(n13933) );
  mux2_1 U21089 ( .ip1(\LUT[29][2] ), .ip2(n17643), .s(n17622), .op(n13932) );
  mux2_1 U21090 ( .ip1(\LUT[29][1] ), .ip2(n17644), .s(n17622), .op(n13931) );
  mux2_1 U21091 ( .ip1(\LUT[29][0] ), .ip2(n17646), .s(n17622), .op(n13930) );
  mux2_1 U21092 ( .ip1(\LUT[28][15] ), .ip2(d[15]), .s(n17623), .op(n13929) );
  mux2_1 U21093 ( .ip1(\LUT[28][14] ), .ip2(d[14]), .s(n17623), .op(n13928) );
  mux2_1 U21094 ( .ip1(\LUT[28][13] ), .ip2(d[13]), .s(n17623), .op(n13927) );
  mux2_1 U21095 ( .ip1(\LUT[28][12] ), .ip2(d[12]), .s(n17623), .op(n13926) );
  mux2_1 U21096 ( .ip1(\LUT[28][11] ), .ip2(d[11]), .s(n17623), .op(n13925) );
  mux2_1 U21097 ( .ip1(\LUT[28][10] ), .ip2(d[10]), .s(n17623), .op(n13924) );
  mux2_1 U21098 ( .ip1(\LUT[28][9] ), .ip2(d[9]), .s(n17623), .op(n13923) );
  mux2_1 U21099 ( .ip1(\LUT[28][8] ), .ip2(d[8]), .s(n17623), .op(n13922) );
  mux2_1 U21100 ( .ip1(\LUT[28][7] ), .ip2(d[7]), .s(n17623), .op(n13921) );
  mux2_1 U21101 ( .ip1(\LUT[28][6] ), .ip2(d[6]), .s(n17623), .op(n13920) );
  mux2_1 U21102 ( .ip1(\LUT[28][5] ), .ip2(d[5]), .s(n17624), .op(n13919) );
  mux2_1 U21103 ( .ip1(\LUT[28][4] ), .ip2(d[4]), .s(n17624), .op(n13918) );
  mux2_1 U21104 ( .ip1(\LUT[28][3] ), .ip2(d[3]), .s(n17624), .op(n13917) );
  mux2_1 U21105 ( .ip1(\LUT[28][2] ), .ip2(d[2]), .s(n17624), .op(n13916) );
  mux2_1 U21106 ( .ip1(\LUT[28][1] ), .ip2(d[1]), .s(n17624), .op(n13915) );
  mux2_1 U21107 ( .ip1(\LUT[28][0] ), .ip2(d[0]), .s(n17624), .op(n13914) );
  mux2_1 U21108 ( .ip1(\LUT[27][15] ), .ip2(n17629), .s(n17625), .op(n13913)
         );
  mux2_1 U21109 ( .ip1(\LUT[27][14] ), .ip2(n17630), .s(n17625), .op(n13912)
         );
  mux2_1 U21110 ( .ip1(\LUT[27][13] ), .ip2(n17631), .s(n17625), .op(n13911)
         );
  mux2_1 U21111 ( .ip1(\LUT[27][12] ), .ip2(n17632), .s(n17625), .op(n13910)
         );
  mux2_1 U21112 ( .ip1(\LUT[27][11] ), .ip2(n17633), .s(n17625), .op(n13909)
         );
  mux2_1 U21113 ( .ip1(\LUT[27][10] ), .ip2(n17634), .s(n17625), .op(n13908)
         );
  mux2_1 U21114 ( .ip1(\LUT[27][9] ), .ip2(n17635), .s(n17625), .op(n13907) );
  mux2_1 U21115 ( .ip1(\LUT[27][8] ), .ip2(n17636), .s(n17625), .op(n13906) );
  mux2_1 U21116 ( .ip1(\LUT[27][7] ), .ip2(n17637), .s(n17625), .op(n13905) );
  mux2_1 U21117 ( .ip1(\LUT[27][6] ), .ip2(n17639), .s(n17625), .op(n13904) );
  mux2_1 U21118 ( .ip1(\LUT[27][5] ), .ip2(n17640), .s(n17626), .op(n13903) );
  mux2_1 U21119 ( .ip1(\LUT[27][4] ), .ip2(n17641), .s(n17626), .op(n13902) );
  mux2_1 U21120 ( .ip1(\LUT[27][3] ), .ip2(n17642), .s(n17626), .op(n13901) );
  mux2_1 U21121 ( .ip1(\LUT[27][2] ), .ip2(n17643), .s(n17626), .op(n13900) );
  mux2_1 U21122 ( .ip1(\LUT[27][1] ), .ip2(n17644), .s(n17626), .op(n13899) );
  mux2_1 U21123 ( .ip1(\LUT[27][0] ), .ip2(n17646), .s(n17626), .op(n13898) );
  mux2_1 U21124 ( .ip1(\LUT[26][15] ), .ip2(d[15]), .s(n17627), .op(n13897) );
  mux2_1 U21125 ( .ip1(\LUT[26][14] ), .ip2(d[14]), .s(n17627), .op(n13896) );
  mux2_1 U21126 ( .ip1(\LUT[26][13] ), .ip2(d[13]), .s(n17627), .op(n13895) );
  mux2_1 U21127 ( .ip1(\LUT[26][12] ), .ip2(d[12]), .s(n17627), .op(n13894) );
  mux2_1 U21128 ( .ip1(\LUT[26][11] ), .ip2(d[11]), .s(n17627), .op(n13893) );
  mux2_1 U21129 ( .ip1(\LUT[26][10] ), .ip2(d[10]), .s(n17627), .op(n13892) );
  mux2_1 U21130 ( .ip1(\LUT[26][9] ), .ip2(d[9]), .s(n17627), .op(n13891) );
  mux2_1 U21131 ( .ip1(\LUT[26][8] ), .ip2(d[8]), .s(n17627), .op(n13890) );
  mux2_1 U21132 ( .ip1(\LUT[26][7] ), .ip2(d[7]), .s(n17627), .op(n13889) );
  mux2_1 U21133 ( .ip1(\LUT[26][6] ), .ip2(d[6]), .s(n17627), .op(n13888) );
  mux2_1 U21134 ( .ip1(\LUT[26][5] ), .ip2(d[5]), .s(n17628), .op(n13887) );
  mux2_1 U21135 ( .ip1(\LUT[26][4] ), .ip2(d[4]), .s(n17628), .op(n13886) );
  mux2_1 U21136 ( .ip1(\LUT[26][3] ), .ip2(d[3]), .s(n17628), .op(n13885) );
  mux2_1 U21137 ( .ip1(\LUT[26][2] ), .ip2(d[2]), .s(n17628), .op(n13884) );
  mux2_1 U21138 ( .ip1(\LUT[26][1] ), .ip2(d[1]), .s(n17628), .op(n13883) );
  mux2_1 U21139 ( .ip1(\LUT[26][0] ), .ip2(d[0]), .s(n17628), .op(n13882) );
  mux2_1 U21140 ( .ip1(\LUT[25][15] ), .ip2(n17629), .s(n17638), .op(n13881)
         );
  mux2_1 U21141 ( .ip1(\LUT[25][14] ), .ip2(n17630), .s(n17638), .op(n13880)
         );
  mux2_1 U21142 ( .ip1(\LUT[25][13] ), .ip2(n17631), .s(n17638), .op(n13879)
         );
  mux2_1 U21143 ( .ip1(\LUT[25][12] ), .ip2(n17632), .s(n17638), .op(n13878)
         );
  mux2_1 U21144 ( .ip1(\LUT[25][11] ), .ip2(n17633), .s(n17638), .op(n13877)
         );
  mux2_1 U21145 ( .ip1(\LUT[25][10] ), .ip2(n17634), .s(n17638), .op(n13876)
         );
  mux2_1 U21146 ( .ip1(\LUT[25][9] ), .ip2(n17635), .s(n17638), .op(n13875) );
  mux2_1 U21147 ( .ip1(\LUT[25][8] ), .ip2(n17636), .s(n17638), .op(n13874) );
  mux2_1 U21148 ( .ip1(\LUT[25][7] ), .ip2(n17637), .s(n17638), .op(n13873) );
  mux2_1 U21149 ( .ip1(\LUT[25][6] ), .ip2(n17639), .s(n17638), .op(n13872) );
  mux2_1 U21150 ( .ip1(\LUT[25][5] ), .ip2(n17640), .s(n17645), .op(n13871) );
  mux2_1 U21151 ( .ip1(\LUT[25][4] ), .ip2(n17641), .s(n17645), .op(n13870) );
  mux2_1 U21152 ( .ip1(\LUT[25][3] ), .ip2(n17642), .s(n17645), .op(n13869) );
  mux2_1 U21153 ( .ip1(\LUT[25][2] ), .ip2(n17643), .s(n17645), .op(n13868) );
  mux2_1 U21154 ( .ip1(\LUT[25][1] ), .ip2(n17644), .s(n17645), .op(n13867) );
  mux2_1 U21155 ( .ip1(\LUT[25][0] ), .ip2(n17646), .s(n17645), .op(n13866) );
  mux2_1 U21156 ( .ip1(\LUT[24][15] ), .ip2(n17629), .s(n17647), .op(n13865)
         );
  mux2_1 U21157 ( .ip1(\LUT[24][14] ), .ip2(n17630), .s(n17647), .op(n13864)
         );
  mux2_1 U21158 ( .ip1(\LUT[24][13] ), .ip2(n17631), .s(n17647), .op(n13863)
         );
  mux2_1 U21159 ( .ip1(\LUT[24][12] ), .ip2(n17632), .s(n17647), .op(n13862)
         );
  mux2_1 U21160 ( .ip1(\LUT[24][11] ), .ip2(n17633), .s(n17647), .op(n13861)
         );
  mux2_1 U21161 ( .ip1(\LUT[24][10] ), .ip2(n17634), .s(n17647), .op(n13860)
         );
  mux2_1 U21162 ( .ip1(\LUT[24][9] ), .ip2(n17635), .s(n17647), .op(n13859) );
  mux2_1 U21163 ( .ip1(\LUT[24][8] ), .ip2(n17636), .s(n17647), .op(n13858) );
  mux2_1 U21164 ( .ip1(\LUT[24][7] ), .ip2(n17637), .s(n17647), .op(n13857) );
  mux2_1 U21165 ( .ip1(\LUT[24][6] ), .ip2(n17639), .s(n17647), .op(n13856) );
  mux2_1 U21166 ( .ip1(\LUT[24][5] ), .ip2(n17640), .s(n17648), .op(n13855) );
  mux2_1 U21167 ( .ip1(\LUT[24][4] ), .ip2(n17641), .s(n17648), .op(n13854) );
  mux2_1 U21168 ( .ip1(\LUT[24][3] ), .ip2(n17642), .s(n17648), .op(n13853) );
  mux2_1 U21169 ( .ip1(\LUT[24][2] ), .ip2(n17643), .s(n17648), .op(n13852) );
  mux2_1 U21170 ( .ip1(\LUT[24][1] ), .ip2(n17644), .s(n17648), .op(n13851) );
  mux2_1 U21171 ( .ip1(\LUT[24][0] ), .ip2(n17646), .s(n17648), .op(n13850) );
  mux2_1 U21172 ( .ip1(\LUT[23][15] ), .ip2(n17629), .s(n17649), .op(n13849)
         );
  mux2_1 U21173 ( .ip1(\LUT[23][14] ), .ip2(n17630), .s(n17649), .op(n13848)
         );
  mux2_1 U21174 ( .ip1(\LUT[23][13] ), .ip2(n17631), .s(n17649), .op(n13847)
         );
  mux2_1 U21175 ( .ip1(\LUT[23][12] ), .ip2(n17632), .s(n17649), .op(n13846)
         );
  mux2_1 U21176 ( .ip1(\LUT[23][11] ), .ip2(n17633), .s(n17649), .op(n13845)
         );
  mux2_1 U21177 ( .ip1(\LUT[23][10] ), .ip2(n17634), .s(n17649), .op(n13844)
         );
  mux2_1 U21178 ( .ip1(\LUT[23][9] ), .ip2(n17635), .s(n17649), .op(n13843) );
  mux2_1 U21179 ( .ip1(\LUT[23][8] ), .ip2(n17636), .s(n17649), .op(n13842) );
  mux2_1 U21180 ( .ip1(\LUT[23][7] ), .ip2(n17637), .s(n17649), .op(n13841) );
  mux2_1 U21181 ( .ip1(\LUT[23][6] ), .ip2(n17639), .s(n17649), .op(n13840) );
  mux2_1 U21182 ( .ip1(\LUT[23][5] ), .ip2(n17640), .s(n17650), .op(n13839) );
  mux2_1 U21183 ( .ip1(\LUT[23][4] ), .ip2(n17641), .s(n17650), .op(n13838) );
  mux2_1 U21184 ( .ip1(\LUT[23][3] ), .ip2(n17642), .s(n17650), .op(n13837) );
  mux2_1 U21185 ( .ip1(\LUT[23][2] ), .ip2(n17643), .s(n17650), .op(n13836) );
  mux2_1 U21186 ( .ip1(\LUT[23][1] ), .ip2(n17644), .s(n17650), .op(n13835) );
  mux2_1 U21187 ( .ip1(\LUT[23][0] ), .ip2(n17646), .s(n17650), .op(n13834) );
  mux2_1 U21188 ( .ip1(\LUT[22][15] ), .ip2(n17629), .s(n17651), .op(n13833)
         );
  mux2_1 U21189 ( .ip1(\LUT[22][14] ), .ip2(n17630), .s(n17651), .op(n13832)
         );
  mux2_1 U21190 ( .ip1(\LUT[22][13] ), .ip2(n17631), .s(n17651), .op(n13831)
         );
  mux2_1 U21191 ( .ip1(\LUT[22][12] ), .ip2(n17632), .s(n17651), .op(n13830)
         );
  mux2_1 U21192 ( .ip1(\LUT[22][11] ), .ip2(n17633), .s(n17651), .op(n13829)
         );
  mux2_1 U21193 ( .ip1(\LUT[22][10] ), .ip2(n17634), .s(n17651), .op(n13828)
         );
  mux2_1 U21194 ( .ip1(\LUT[22][9] ), .ip2(n17635), .s(n17651), .op(n13827) );
  mux2_1 U21195 ( .ip1(\LUT[22][8] ), .ip2(n17636), .s(n17651), .op(n13826) );
  mux2_1 U21196 ( .ip1(\LUT[22][7] ), .ip2(n17637), .s(n17651), .op(n13825) );
  mux2_1 U21197 ( .ip1(\LUT[22][6] ), .ip2(n17639), .s(n17651), .op(n13824) );
  mux2_1 U21198 ( .ip1(\LUT[22][5] ), .ip2(n17640), .s(n17652), .op(n13823) );
  mux2_1 U21199 ( .ip1(\LUT[22][4] ), .ip2(n17641), .s(n17652), .op(n13822) );
  mux2_1 U21200 ( .ip1(\LUT[22][3] ), .ip2(n17642), .s(n17652), .op(n13821) );
  mux2_1 U21201 ( .ip1(\LUT[22][2] ), .ip2(n17643), .s(n17652), .op(n13820) );
  mux2_1 U21202 ( .ip1(\LUT[22][1] ), .ip2(n17644), .s(n17652), .op(n13819) );
  mux2_1 U21203 ( .ip1(\LUT[22][0] ), .ip2(n17646), .s(n17652), .op(n13818) );
  mux2_1 U21204 ( .ip1(\LUT[21][15] ), .ip2(n17629), .s(n17653), .op(n13817)
         );
  mux2_1 U21205 ( .ip1(\LUT[21][14] ), .ip2(n17630), .s(n17653), .op(n13816)
         );
  mux2_1 U21206 ( .ip1(\LUT[21][13] ), .ip2(n17631), .s(n17653), .op(n13815)
         );
  mux2_1 U21207 ( .ip1(\LUT[21][12] ), .ip2(n17632), .s(n17653), .op(n13814)
         );
  mux2_1 U21208 ( .ip1(\LUT[21][11] ), .ip2(n17633), .s(n17653), .op(n13813)
         );
  mux2_1 U21209 ( .ip1(\LUT[21][10] ), .ip2(n17634), .s(n17653), .op(n13812)
         );
  mux2_1 U21210 ( .ip1(\LUT[21][9] ), .ip2(n17635), .s(n17653), .op(n13811) );
  mux2_1 U21211 ( .ip1(\LUT[21][8] ), .ip2(n17636), .s(n17653), .op(n13810) );
  mux2_1 U21212 ( .ip1(\LUT[21][7] ), .ip2(n17637), .s(n17653), .op(n13809) );
  mux2_1 U21213 ( .ip1(\LUT[21][6] ), .ip2(n17639), .s(n17653), .op(n13808) );
  mux2_1 U21214 ( .ip1(\LUT[21][5] ), .ip2(n17640), .s(n17654), .op(n13807) );
  mux2_1 U21215 ( .ip1(\LUT[21][4] ), .ip2(n17641), .s(n17654), .op(n13806) );
  mux2_1 U21216 ( .ip1(\LUT[21][3] ), .ip2(n17642), .s(n17654), .op(n13805) );
  mux2_1 U21217 ( .ip1(\LUT[21][2] ), .ip2(n17643), .s(n17654), .op(n13804) );
  mux2_1 U21218 ( .ip1(\LUT[21][1] ), .ip2(n17644), .s(n17654), .op(n13803) );
  mux2_1 U21219 ( .ip1(\LUT[21][0] ), .ip2(n17646), .s(n17654), .op(n13802) );
  mux2_1 U21220 ( .ip1(\LUT[20][15] ), .ip2(n17629), .s(n17655), .op(n13801)
         );
  mux2_1 U21221 ( .ip1(\LUT[20][14] ), .ip2(n17630), .s(n17655), .op(n13800)
         );
  mux2_1 U21222 ( .ip1(\LUT[20][13] ), .ip2(n17631), .s(n17655), .op(n13799)
         );
  mux2_1 U21223 ( .ip1(\LUT[20][12] ), .ip2(n17632), .s(n17655), .op(n13798)
         );
  mux2_1 U21224 ( .ip1(\LUT[20][11] ), .ip2(n17633), .s(n17655), .op(n13797)
         );
  mux2_1 U21225 ( .ip1(\LUT[20][10] ), .ip2(n17634), .s(n17655), .op(n13796)
         );
  mux2_1 U21226 ( .ip1(\LUT[20][9] ), .ip2(n17635), .s(n17655), .op(n13795) );
  mux2_1 U21227 ( .ip1(\LUT[20][8] ), .ip2(n17636), .s(n17655), .op(n13794) );
  mux2_1 U21228 ( .ip1(\LUT[20][7] ), .ip2(n17637), .s(n17655), .op(n13793) );
  mux2_1 U21229 ( .ip1(\LUT[20][6] ), .ip2(n17639), .s(n17655), .op(n13792) );
  mux2_1 U21230 ( .ip1(\LUT[20][5] ), .ip2(n17640), .s(n17656), .op(n13791) );
  mux2_1 U21231 ( .ip1(\LUT[20][4] ), .ip2(n17641), .s(n17656), .op(n13790) );
  mux2_1 U21232 ( .ip1(\LUT[20][3] ), .ip2(n17642), .s(n17656), .op(n13789) );
  mux2_1 U21233 ( .ip1(\LUT[20][2] ), .ip2(n17643), .s(n17656), .op(n13788) );
  mux2_1 U21234 ( .ip1(\LUT[20][1] ), .ip2(n17644), .s(n17656), .op(n13787) );
  mux2_1 U21235 ( .ip1(\LUT[20][0] ), .ip2(n17646), .s(n17656), .op(n13786) );
  mux2_1 U21236 ( .ip1(\LUT[19][15] ), .ip2(n17541), .s(n17657), .op(n13785)
         );
  mux2_1 U21237 ( .ip1(\LUT[19][14] ), .ip2(n17542), .s(n17657), .op(n13784)
         );
  mux2_1 U21238 ( .ip1(\LUT[19][13] ), .ip2(n17543), .s(n17657), .op(n13783)
         );
  mux2_1 U21239 ( .ip1(\LUT[19][12] ), .ip2(n17544), .s(n17657), .op(n13782)
         );
  mux2_1 U21240 ( .ip1(\LUT[19][11] ), .ip2(n17545), .s(n17657), .op(n13781)
         );
  mux2_1 U21241 ( .ip1(\LUT[19][10] ), .ip2(n17546), .s(n17657), .op(n13780)
         );
  mux2_1 U21242 ( .ip1(\LUT[19][9] ), .ip2(n17547), .s(n17657), .op(n13779) );
  mux2_1 U21243 ( .ip1(\LUT[19][8] ), .ip2(n17548), .s(n17657), .op(n13778) );
  mux2_1 U21244 ( .ip1(\LUT[19][7] ), .ip2(n17549), .s(n17657), .op(n13777) );
  mux2_1 U21245 ( .ip1(\LUT[19][6] ), .ip2(n17551), .s(n17657), .op(n13776) );
  mux2_1 U21246 ( .ip1(\LUT[19][5] ), .ip2(n17552), .s(n17658), .op(n13775) );
  mux2_1 U21247 ( .ip1(\LUT[19][4] ), .ip2(n17553), .s(n17658), .op(n13774) );
  mux2_1 U21248 ( .ip1(\LUT[19][3] ), .ip2(n17554), .s(n17658), .op(n13773) );
  mux2_1 U21249 ( .ip1(\LUT[19][2] ), .ip2(n17555), .s(n17658), .op(n13772) );
  mux2_1 U21250 ( .ip1(\LUT[19][1] ), .ip2(n17556), .s(n17658), .op(n13771) );
  mux2_1 U21251 ( .ip1(\LUT[19][0] ), .ip2(n17558), .s(n17658), .op(n13770) );
  mux2_1 U21252 ( .ip1(\LUT[18][15] ), .ip2(d[15]), .s(n17659), .op(n13769) );
  mux2_1 U21253 ( .ip1(\LUT[18][14] ), .ip2(d[14]), .s(n17659), .op(n13768) );
  mux2_1 U21254 ( .ip1(\LUT[18][13] ), .ip2(d[13]), .s(n17659), .op(n13767) );
  mux2_1 U21255 ( .ip1(\LUT[18][12] ), .ip2(d[12]), .s(n17659), .op(n13766) );
  mux2_1 U21256 ( .ip1(\LUT[18][11] ), .ip2(d[11]), .s(n17659), .op(n13765) );
  mux2_1 U21257 ( .ip1(\LUT[18][10] ), .ip2(d[10]), .s(n17659), .op(n13764) );
  mux2_1 U21258 ( .ip1(\LUT[18][9] ), .ip2(d[9]), .s(n17659), .op(n13763) );
  mux2_1 U21259 ( .ip1(\LUT[18][8] ), .ip2(d[8]), .s(n17659), .op(n13762) );
  mux2_1 U21260 ( .ip1(\LUT[18][7] ), .ip2(d[7]), .s(n17659), .op(n13761) );
  mux2_1 U21261 ( .ip1(\LUT[18][6] ), .ip2(d[6]), .s(n17659), .op(n13760) );
  mux2_1 U21262 ( .ip1(\LUT[18][5] ), .ip2(d[5]), .s(n17660), .op(n13759) );
  mux2_1 U21263 ( .ip1(\LUT[18][4] ), .ip2(d[4]), .s(n17660), .op(n13758) );
  mux2_1 U21264 ( .ip1(\LUT[18][3] ), .ip2(d[3]), .s(n17660), .op(n13757) );
  mux2_1 U21265 ( .ip1(\LUT[18][2] ), .ip2(d[2]), .s(n17660), .op(n13756) );
  mux2_1 U21266 ( .ip1(\LUT[18][1] ), .ip2(d[1]), .s(n17660), .op(n13755) );
  mux2_1 U21267 ( .ip1(\LUT[18][0] ), .ip2(d[0]), .s(n17660), .op(n13754) );
  mux2_1 U21268 ( .ip1(\LUT[17][15] ), .ip2(n17629), .s(n17661), .op(n13753)
         );
  mux2_1 U21269 ( .ip1(\LUT[17][14] ), .ip2(n17630), .s(n17661), .op(n13752)
         );
  mux2_1 U21270 ( .ip1(\LUT[17][13] ), .ip2(n17631), .s(n17661), .op(n13751)
         );
  mux2_1 U21271 ( .ip1(\LUT[17][12] ), .ip2(n17632), .s(n17661), .op(n13750)
         );
  mux2_1 U21272 ( .ip1(\LUT[17][11] ), .ip2(n17633), .s(n17661), .op(n13749)
         );
  mux2_1 U21273 ( .ip1(\LUT[17][10] ), .ip2(n17634), .s(n17661), .op(n13748)
         );
  mux2_1 U21274 ( .ip1(\LUT[17][9] ), .ip2(n17635), .s(n17661), .op(n13747) );
  mux2_1 U21275 ( .ip1(\LUT[17][8] ), .ip2(n17636), .s(n17661), .op(n13746) );
  mux2_1 U21276 ( .ip1(\LUT[17][7] ), .ip2(n17637), .s(n17661), .op(n13745) );
  mux2_1 U21277 ( .ip1(\LUT[17][6] ), .ip2(n17639), .s(n17661), .op(n13744) );
  mux2_1 U21278 ( .ip1(\LUT[17][5] ), .ip2(n17640), .s(n17662), .op(n13743) );
  mux2_1 U21279 ( .ip1(\LUT[17][4] ), .ip2(n17641), .s(n17662), .op(n13742) );
  mux2_1 U21280 ( .ip1(\LUT[17][3] ), .ip2(n17642), .s(n17662), .op(n13741) );
  mux2_1 U21281 ( .ip1(\LUT[17][2] ), .ip2(n17643), .s(n17662), .op(n13740) );
  mux2_1 U21282 ( .ip1(\LUT[17][1] ), .ip2(n17644), .s(n17662), .op(n13739) );
  mux2_1 U21283 ( .ip1(\LUT[17][0] ), .ip2(n17646), .s(n17662), .op(n13738) );
  mux2_1 U21284 ( .ip1(\LUT[16][15] ), .ip2(d[15]), .s(n17663), .op(n13737) );
  mux2_1 U21285 ( .ip1(\LUT[16][14] ), .ip2(d[14]), .s(n17663), .op(n13736) );
  mux2_1 U21286 ( .ip1(\LUT[16][13] ), .ip2(d[13]), .s(n17663), .op(n13735) );
  mux2_1 U21287 ( .ip1(\LUT[16][12] ), .ip2(d[12]), .s(n17663), .op(n13734) );
  mux2_1 U21288 ( .ip1(\LUT[16][11] ), .ip2(d[11]), .s(n17663), .op(n13733) );
  mux2_1 U21289 ( .ip1(\LUT[16][10] ), .ip2(d[10]), .s(n17663), .op(n13732) );
  mux2_1 U21290 ( .ip1(\LUT[16][9] ), .ip2(d[9]), .s(n17663), .op(n13731) );
  mux2_1 U21291 ( .ip1(\LUT[16][8] ), .ip2(d[8]), .s(n17663), .op(n13730) );
  mux2_1 U21292 ( .ip1(\LUT[16][7] ), .ip2(d[7]), .s(n17663), .op(n13729) );
  mux2_1 U21293 ( .ip1(\LUT[16][6] ), .ip2(d[6]), .s(n17663), .op(n13728) );
  mux2_1 U21294 ( .ip1(\LUT[16][5] ), .ip2(d[5]), .s(n17664), .op(n13727) );
  mux2_1 U21295 ( .ip1(\LUT[16][4] ), .ip2(d[4]), .s(n17664), .op(n13726) );
  mux2_1 U21296 ( .ip1(\LUT[16][3] ), .ip2(d[3]), .s(n17664), .op(n13725) );
  mux2_1 U21297 ( .ip1(\LUT[16][2] ), .ip2(d[2]), .s(n17664), .op(n13724) );
  mux2_1 U21298 ( .ip1(\LUT[16][1] ), .ip2(d[1]), .s(n17664), .op(n13723) );
  mux2_1 U21299 ( .ip1(\LUT[16][0] ), .ip2(d[0]), .s(n17664), .op(n13722) );
  mux2_1 U21300 ( .ip1(\LUT[15][15] ), .ip2(d[15]), .s(n17665), .op(n13721) );
  mux2_1 U21301 ( .ip1(\LUT[15][14] ), .ip2(d[14]), .s(n17665), .op(n13720) );
  mux2_1 U21302 ( .ip1(\LUT[15][13] ), .ip2(d[13]), .s(n17665), .op(n13719) );
  mux2_1 U21303 ( .ip1(\LUT[15][12] ), .ip2(d[12]), .s(n17665), .op(n13718) );
  mux2_1 U21304 ( .ip1(\LUT[15][11] ), .ip2(d[11]), .s(n17665), .op(n13717) );
  mux2_1 U21305 ( .ip1(\LUT[15][10] ), .ip2(d[10]), .s(n17665), .op(n13716) );
  mux2_1 U21306 ( .ip1(\LUT[15][9] ), .ip2(d[9]), .s(n17665), .op(n13715) );
  mux2_1 U21307 ( .ip1(\LUT[15][8] ), .ip2(d[8]), .s(n17665), .op(n13714) );
  mux2_1 U21308 ( .ip1(\LUT[15][7] ), .ip2(d[7]), .s(n17665), .op(n13713) );
  mux2_1 U21309 ( .ip1(\LUT[15][6] ), .ip2(d[6]), .s(n17665), .op(n13712) );
  mux2_1 U21310 ( .ip1(\LUT[15][5] ), .ip2(d[5]), .s(n17666), .op(n13711) );
  mux2_1 U21311 ( .ip1(\LUT[15][4] ), .ip2(d[4]), .s(n17666), .op(n13710) );
  mux2_1 U21312 ( .ip1(\LUT[15][3] ), .ip2(d[3]), .s(n17666), .op(n13709) );
  mux2_1 U21313 ( .ip1(\LUT[15][2] ), .ip2(d[2]), .s(n17666), .op(n13708) );
  mux2_1 U21314 ( .ip1(\LUT[15][1] ), .ip2(d[1]), .s(n17666), .op(n13707) );
  mux2_1 U21315 ( .ip1(\LUT[15][0] ), .ip2(d[0]), .s(n17666), .op(n13706) );
  mux2_1 U21316 ( .ip1(\LUT[14][15] ), .ip2(n17541), .s(n17667), .op(n13705)
         );
  mux2_1 U21317 ( .ip1(\LUT[14][14] ), .ip2(n17542), .s(n17667), .op(n13704)
         );
  mux2_1 U21318 ( .ip1(\LUT[14][13] ), .ip2(n17543), .s(n17667), .op(n13703)
         );
  mux2_1 U21319 ( .ip1(\LUT[14][12] ), .ip2(n17544), .s(n17667), .op(n13702)
         );
  mux2_1 U21320 ( .ip1(\LUT[14][11] ), .ip2(n17545), .s(n17667), .op(n13701)
         );
  mux2_1 U21321 ( .ip1(\LUT[14][10] ), .ip2(n17546), .s(n17667), .op(n13700)
         );
  mux2_1 U21322 ( .ip1(\LUT[14][9] ), .ip2(n17547), .s(n17667), .op(n13699) );
  mux2_1 U21323 ( .ip1(\LUT[14][8] ), .ip2(n17548), .s(n17667), .op(n13698) );
  mux2_1 U21324 ( .ip1(\LUT[14][7] ), .ip2(n17549), .s(n17667), .op(n13697) );
  mux2_1 U21325 ( .ip1(\LUT[14][6] ), .ip2(n17551), .s(n17667), .op(n13696) );
  mux2_1 U21326 ( .ip1(\LUT[14][5] ), .ip2(n17552), .s(n17668), .op(n13695) );
  mux2_1 U21327 ( .ip1(\LUT[14][4] ), .ip2(n17553), .s(n17668), .op(n13694) );
  mux2_1 U21328 ( .ip1(\LUT[14][3] ), .ip2(n17554), .s(n17668), .op(n13693) );
  mux2_1 U21329 ( .ip1(\LUT[14][2] ), .ip2(n17555), .s(n17668), .op(n13692) );
  mux2_1 U21330 ( .ip1(\LUT[14][1] ), .ip2(n17556), .s(n17668), .op(n13691) );
  mux2_1 U21331 ( .ip1(\LUT[14][0] ), .ip2(n17558), .s(n17668), .op(n13690) );
  mux2_1 U21332 ( .ip1(\LUT[13][15] ), .ip2(n17629), .s(n17669), .op(n13689)
         );
  mux2_1 U21333 ( .ip1(\LUT[13][14] ), .ip2(n17630), .s(n17669), .op(n13688)
         );
  mux2_1 U21334 ( .ip1(\LUT[13][13] ), .ip2(n17631), .s(n17669), .op(n13687)
         );
  mux2_1 U21335 ( .ip1(\LUT[13][12] ), .ip2(n17632), .s(n17669), .op(n13686)
         );
  mux2_1 U21336 ( .ip1(\LUT[13][11] ), .ip2(n17633), .s(n17669), .op(n13685)
         );
  mux2_1 U21337 ( .ip1(\LUT[13][10] ), .ip2(n17634), .s(n17669), .op(n13684)
         );
  mux2_1 U21338 ( .ip1(\LUT[13][9] ), .ip2(n17635), .s(n17669), .op(n13683) );
  mux2_1 U21339 ( .ip1(\LUT[13][8] ), .ip2(n17636), .s(n17669), .op(n13682) );
  mux2_1 U21340 ( .ip1(\LUT[13][7] ), .ip2(n17637), .s(n17669), .op(n13681) );
  mux2_1 U21341 ( .ip1(\LUT[13][6] ), .ip2(n17639), .s(n17669), .op(n13680) );
  mux2_1 U21342 ( .ip1(\LUT[13][5] ), .ip2(n17640), .s(n17670), .op(n13679) );
  mux2_1 U21343 ( .ip1(\LUT[13][4] ), .ip2(n17641), .s(n17670), .op(n13678) );
  mux2_1 U21344 ( .ip1(\LUT[13][3] ), .ip2(n17642), .s(n17670), .op(n13677) );
  mux2_1 U21345 ( .ip1(\LUT[13][2] ), .ip2(n17643), .s(n17670), .op(n13676) );
  mux2_1 U21346 ( .ip1(\LUT[13][1] ), .ip2(n17644), .s(n17670), .op(n13675) );
  mux2_1 U21347 ( .ip1(\LUT[13][0] ), .ip2(n17646), .s(n17670), .op(n13674) );
  mux2_1 U21348 ( .ip1(\LUT[12][15] ), .ip2(d[15]), .s(n17671), .op(n13673) );
  mux2_1 U21349 ( .ip1(\LUT[12][14] ), .ip2(d[14]), .s(n17671), .op(n13672) );
  mux2_1 U21350 ( .ip1(\LUT[12][13] ), .ip2(d[13]), .s(n17671), .op(n13671) );
  mux2_1 U21351 ( .ip1(\LUT[12][12] ), .ip2(d[12]), .s(n17671), .op(n13670) );
  mux2_1 U21352 ( .ip1(\LUT[12][11] ), .ip2(d[11]), .s(n17671), .op(n13669) );
  mux2_1 U21353 ( .ip1(\LUT[12][10] ), .ip2(d[10]), .s(n17671), .op(n13668) );
  mux2_1 U21354 ( .ip1(\LUT[12][9] ), .ip2(d[9]), .s(n17671), .op(n13667) );
  mux2_1 U21355 ( .ip1(\LUT[12][8] ), .ip2(d[8]), .s(n17671), .op(n13666) );
  mux2_1 U21356 ( .ip1(\LUT[12][7] ), .ip2(d[7]), .s(n17671), .op(n13665) );
  mux2_1 U21357 ( .ip1(\LUT[12][6] ), .ip2(d[6]), .s(n17671), .op(n13664) );
  mux2_1 U21358 ( .ip1(\LUT[12][5] ), .ip2(d[5]), .s(n17672), .op(n13663) );
  mux2_1 U21359 ( .ip1(\LUT[12][4] ), .ip2(d[4]), .s(n17672), .op(n13662) );
  mux2_1 U21360 ( .ip1(\LUT[12][3] ), .ip2(d[3]), .s(n17672), .op(n13661) );
  mux2_1 U21361 ( .ip1(\LUT[12][2] ), .ip2(d[2]), .s(n17672), .op(n13660) );
  mux2_1 U21362 ( .ip1(\LUT[12][1] ), .ip2(d[1]), .s(n17672), .op(n13659) );
  mux2_1 U21363 ( .ip1(\LUT[12][0] ), .ip2(d[0]), .s(n17672), .op(n13658) );
  mux2_1 U21364 ( .ip1(\LUT[11][15] ), .ip2(n17451), .s(n17673), .op(n13657)
         );
  mux2_1 U21365 ( .ip1(\LUT[11][14] ), .ip2(n17452), .s(n17673), .op(n13656)
         );
  mux2_1 U21366 ( .ip1(\LUT[11][13] ), .ip2(n17453), .s(n17673), .op(n13655)
         );
  mux2_1 U21367 ( .ip1(\LUT[11][12] ), .ip2(n17454), .s(n17673), .op(n13654)
         );
  mux2_1 U21368 ( .ip1(\LUT[11][11] ), .ip2(n17455), .s(n17673), .op(n13653)
         );
  mux2_1 U21369 ( .ip1(\LUT[11][10] ), .ip2(n17456), .s(n17673), .op(n13652)
         );
  mux2_1 U21370 ( .ip1(\LUT[11][9] ), .ip2(n17457), .s(n17673), .op(n13651) );
  mux2_1 U21371 ( .ip1(\LUT[11][8] ), .ip2(n17458), .s(n17673), .op(n13650) );
  mux2_1 U21372 ( .ip1(\LUT[11][7] ), .ip2(n17459), .s(n17673), .op(n13649) );
  mux2_1 U21373 ( .ip1(\LUT[11][6] ), .ip2(n17461), .s(n17673), .op(n13648) );
  mux2_1 U21374 ( .ip1(\LUT[11][5] ), .ip2(n17462), .s(n17674), .op(n13647) );
  mux2_1 U21375 ( .ip1(\LUT[11][4] ), .ip2(n17463), .s(n17674), .op(n13646) );
  mux2_1 U21376 ( .ip1(\LUT[11][3] ), .ip2(n17464), .s(n17674), .op(n13645) );
  mux2_1 U21377 ( .ip1(\LUT[11][2] ), .ip2(n17465), .s(n17674), .op(n13644) );
  mux2_1 U21378 ( .ip1(\LUT[11][1] ), .ip2(n17466), .s(n17674), .op(n13643) );
  mux2_1 U21379 ( .ip1(\LUT[11][0] ), .ip2(n17468), .s(n17674), .op(n13642) );
  mux2_1 U21380 ( .ip1(\LUT[10][15] ), .ip2(d[15]), .s(n17675), .op(n13641) );
  mux2_1 U21381 ( .ip1(\LUT[10][14] ), .ip2(d[14]), .s(n17675), .op(n13640) );
  mux2_1 U21382 ( .ip1(\LUT[10][13] ), .ip2(d[13]), .s(n17675), .op(n13639) );
  mux2_1 U21383 ( .ip1(\LUT[10][12] ), .ip2(d[12]), .s(n17675), .op(n13638) );
  mux2_1 U21384 ( .ip1(\LUT[10][11] ), .ip2(d[11]), .s(n17675), .op(n13637) );
  mux2_1 U21385 ( .ip1(\LUT[10][10] ), .ip2(d[10]), .s(n17675), .op(n13636) );
  mux2_1 U21386 ( .ip1(\LUT[10][9] ), .ip2(d[9]), .s(n17675), .op(n13635) );
  mux2_1 U21387 ( .ip1(\LUT[10][8] ), .ip2(d[8]), .s(n17675), .op(n13634) );
  mux2_1 U21388 ( .ip1(\LUT[10][7] ), .ip2(d[7]), .s(n17675), .op(n13633) );
  mux2_1 U21389 ( .ip1(\LUT[10][6] ), .ip2(d[6]), .s(n17675), .op(n13632) );
  mux2_1 U21390 ( .ip1(\LUT[10][5] ), .ip2(d[5]), .s(n17676), .op(n13631) );
  mux2_1 U21391 ( .ip1(\LUT[10][4] ), .ip2(d[4]), .s(n17676), .op(n13630) );
  mux2_1 U21392 ( .ip1(\LUT[10][3] ), .ip2(d[3]), .s(n17676), .op(n13629) );
  mux2_1 U21393 ( .ip1(\LUT[10][2] ), .ip2(d[2]), .s(n17676), .op(n13628) );
  mux2_1 U21394 ( .ip1(\LUT[10][1] ), .ip2(d[1]), .s(n17676), .op(n13627) );
  mux2_1 U21395 ( .ip1(\LUT[10][0] ), .ip2(d[0]), .s(n17676), .op(n13626) );
  mux2_1 U21396 ( .ip1(\LUT[9][15] ), .ip2(n17541), .s(n17677), .op(n13625) );
  mux2_1 U21397 ( .ip1(\LUT[9][14] ), .ip2(n17542), .s(n17677), .op(n13624) );
  mux2_1 U21398 ( .ip1(\LUT[9][13] ), .ip2(n17543), .s(n17677), .op(n13623) );
  mux2_1 U21399 ( .ip1(\LUT[9][12] ), .ip2(n17544), .s(n17677), .op(n13622) );
  mux2_1 U21400 ( .ip1(\LUT[9][11] ), .ip2(n17545), .s(n17677), .op(n13621) );
  mux2_1 U21401 ( .ip1(\LUT[9][10] ), .ip2(n17546), .s(n17677), .op(n13620) );
  mux2_1 U21402 ( .ip1(\LUT[9][9] ), .ip2(n17547), .s(n17677), .op(n13619) );
  mux2_1 U21403 ( .ip1(\LUT[9][8] ), .ip2(n17548), .s(n17677), .op(n13618) );
  mux2_1 U21404 ( .ip1(\LUT[9][7] ), .ip2(n17549), .s(n17677), .op(n13617) );
  mux2_1 U21405 ( .ip1(\LUT[9][6] ), .ip2(n17551), .s(n17677), .op(n13616) );
  mux2_1 U21406 ( .ip1(\LUT[9][5] ), .ip2(n17552), .s(n17678), .op(n13615) );
  mux2_1 U21407 ( .ip1(\LUT[9][4] ), .ip2(n17553), .s(n17678), .op(n13614) );
  mux2_1 U21408 ( .ip1(\LUT[9][3] ), .ip2(n17554), .s(n17678), .op(n13613) );
  mux2_1 U21409 ( .ip1(\LUT[9][2] ), .ip2(n17555), .s(n17678), .op(n13612) );
  mux2_1 U21410 ( .ip1(\LUT[9][1] ), .ip2(n17556), .s(n17678), .op(n13611) );
  mux2_1 U21411 ( .ip1(\LUT[9][0] ), .ip2(n17558), .s(n17678), .op(n13610) );
  mux2_1 U21412 ( .ip1(\LUT[8][15] ), .ip2(n17629), .s(n17679), .op(n13609) );
  mux2_1 U21413 ( .ip1(\LUT[8][14] ), .ip2(n17630), .s(n17679), .op(n13608) );
  mux2_1 U21414 ( .ip1(\LUT[8][13] ), .ip2(n17631), .s(n17679), .op(n13607) );
  mux2_1 U21415 ( .ip1(\LUT[8][12] ), .ip2(n17632), .s(n17679), .op(n13606) );
  mux2_1 U21416 ( .ip1(\LUT[8][11] ), .ip2(n17633), .s(n17679), .op(n13605) );
  mux2_1 U21417 ( .ip1(\LUT[8][10] ), .ip2(n17634), .s(n17679), .op(n13604) );
  mux2_1 U21418 ( .ip1(\LUT[8][9] ), .ip2(n17635), .s(n17679), .op(n13603) );
  mux2_1 U21419 ( .ip1(\LUT[8][8] ), .ip2(n17636), .s(n17679), .op(n13602) );
  mux2_1 U21420 ( .ip1(\LUT[8][7] ), .ip2(n17637), .s(n17679), .op(n13601) );
  mux2_1 U21421 ( .ip1(\LUT[8][6] ), .ip2(n17639), .s(n17679), .op(n13600) );
  mux2_1 U21422 ( .ip1(\LUT[8][5] ), .ip2(n17640), .s(n17680), .op(n13599) );
  mux2_1 U21423 ( .ip1(\LUT[8][4] ), .ip2(n17641), .s(n17680), .op(n13598) );
  mux2_1 U21424 ( .ip1(\LUT[8][3] ), .ip2(n17642), .s(n17680), .op(n13597) );
  mux2_1 U21425 ( .ip1(\LUT[8][2] ), .ip2(n17643), .s(n17680), .op(n13596) );
  mux2_1 U21426 ( .ip1(\LUT[8][1] ), .ip2(n17644), .s(n17680), .op(n13595) );
  mux2_1 U21427 ( .ip1(\LUT[8][0] ), .ip2(n17646), .s(n17680), .op(n13594) );
  mux2_1 U21428 ( .ip1(\LUT[7][15] ), .ip2(d[15]), .s(n17681), .op(n13593) );
  mux2_1 U21429 ( .ip1(\LUT[7][14] ), .ip2(d[14]), .s(n17681), .op(n13592) );
  mux2_1 U21430 ( .ip1(\LUT[7][13] ), .ip2(d[13]), .s(n17681), .op(n13591) );
  mux2_1 U21431 ( .ip1(\LUT[7][12] ), .ip2(d[12]), .s(n17681), .op(n13590) );
  mux2_1 U21432 ( .ip1(\LUT[7][11] ), .ip2(d[11]), .s(n17681), .op(n13589) );
  mux2_1 U21433 ( .ip1(\LUT[7][10] ), .ip2(d[10]), .s(n17681), .op(n13588) );
  mux2_1 U21434 ( .ip1(\LUT[7][9] ), .ip2(d[9]), .s(n17681), .op(n13587) );
  mux2_1 U21435 ( .ip1(\LUT[7][8] ), .ip2(d[8]), .s(n17681), .op(n13586) );
  mux2_1 U21436 ( .ip1(\LUT[7][7] ), .ip2(d[7]), .s(n17681), .op(n13585) );
  mux2_1 U21437 ( .ip1(\LUT[7][6] ), .ip2(d[6]), .s(n17681), .op(n13584) );
  mux2_1 U21438 ( .ip1(\LUT[7][5] ), .ip2(d[5]), .s(n17682), .op(n13583) );
  mux2_1 U21439 ( .ip1(\LUT[7][4] ), .ip2(d[4]), .s(n17682), .op(n13582) );
  mux2_1 U21440 ( .ip1(\LUT[7][3] ), .ip2(d[3]), .s(n17682), .op(n13581) );
  mux2_1 U21441 ( .ip1(\LUT[7][2] ), .ip2(d[2]), .s(n17682), .op(n13580) );
  mux2_1 U21442 ( .ip1(\LUT[7][1] ), .ip2(d[1]), .s(n17682), .op(n13579) );
  mux2_1 U21443 ( .ip1(\LUT[7][0] ), .ip2(d[0]), .s(n17682), .op(n13578) );
  mux2_1 U21444 ( .ip1(\LUT[6][15] ), .ip2(n17451), .s(n17683), .op(n13577) );
  mux2_1 U21445 ( .ip1(\LUT[6][14] ), .ip2(n17452), .s(n17683), .op(n13576) );
  mux2_1 U21446 ( .ip1(\LUT[6][13] ), .ip2(n17453), .s(n17683), .op(n13575) );
  mux2_1 U21447 ( .ip1(\LUT[6][12] ), .ip2(n17454), .s(n17683), .op(n13574) );
  mux2_1 U21448 ( .ip1(\LUT[6][11] ), .ip2(n17455), .s(n17683), .op(n13573) );
  mux2_1 U21449 ( .ip1(\LUT[6][10] ), .ip2(n17456), .s(n17683), .op(n13572) );
  mux2_1 U21450 ( .ip1(\LUT[6][9] ), .ip2(n17457), .s(n17683), .op(n13571) );
  mux2_1 U21451 ( .ip1(\LUT[6][8] ), .ip2(n17458), .s(n17683), .op(n13570) );
  mux2_1 U21452 ( .ip1(\LUT[6][7] ), .ip2(n17459), .s(n17683), .op(n13569) );
  mux2_1 U21453 ( .ip1(\LUT[6][6] ), .ip2(n17461), .s(n17683), .op(n13568) );
  mux2_1 U21454 ( .ip1(\LUT[6][5] ), .ip2(n17462), .s(n17684), .op(n13567) );
  mux2_1 U21455 ( .ip1(\LUT[6][4] ), .ip2(n17463), .s(n17684), .op(n13566) );
  mux2_1 U21456 ( .ip1(\LUT[6][3] ), .ip2(n17464), .s(n17684), .op(n13565) );
  mux2_1 U21457 ( .ip1(\LUT[6][2] ), .ip2(n17465), .s(n17684), .op(n13564) );
  mux2_1 U21458 ( .ip1(\LUT[6][1] ), .ip2(n17466), .s(n17684), .op(n13563) );
  mux2_1 U21459 ( .ip1(\LUT[6][0] ), .ip2(n17468), .s(n17684), .op(n13562) );
  mux2_1 U21460 ( .ip1(\LUT[5][15] ), .ip2(n17541), .s(n17685), .op(n13561) );
  mux2_1 U21461 ( .ip1(\LUT[5][14] ), .ip2(n17542), .s(n17685), .op(n13560) );
  mux2_1 U21462 ( .ip1(\LUT[5][13] ), .ip2(n17543), .s(n17685), .op(n13559) );
  mux2_1 U21463 ( .ip1(\LUT[5][12] ), .ip2(n17544), .s(n17685), .op(n13558) );
  mux2_1 U21464 ( .ip1(\LUT[5][11] ), .ip2(n17545), .s(n17685), .op(n13557) );
  mux2_1 U21465 ( .ip1(\LUT[5][10] ), .ip2(n17546), .s(n17685), .op(n13556) );
  mux2_1 U21466 ( .ip1(\LUT[5][9] ), .ip2(n17547), .s(n17685), .op(n13555) );
  mux2_1 U21467 ( .ip1(\LUT[5][8] ), .ip2(n17548), .s(n17685), .op(n13554) );
  mux2_1 U21468 ( .ip1(\LUT[5][7] ), .ip2(n17549), .s(n17685), .op(n13553) );
  mux2_1 U21469 ( .ip1(\LUT[5][6] ), .ip2(n17551), .s(n17685), .op(n13552) );
  mux2_1 U21470 ( .ip1(\LUT[5][5] ), .ip2(n17552), .s(n17686), .op(n13551) );
  mux2_1 U21471 ( .ip1(\LUT[5][4] ), .ip2(n17553), .s(n17686), .op(n13550) );
  mux2_1 U21472 ( .ip1(\LUT[5][3] ), .ip2(n17554), .s(n17686), .op(n13549) );
  mux2_1 U21473 ( .ip1(\LUT[5][2] ), .ip2(n17555), .s(n17686), .op(n13548) );
  mux2_1 U21474 ( .ip1(\LUT[5][1] ), .ip2(n17556), .s(n17686), .op(n13547) );
  mux2_1 U21475 ( .ip1(\LUT[5][0] ), .ip2(n17558), .s(n17686), .op(n13546) );
  mux2_1 U21476 ( .ip1(\LUT[4][15] ), .ip2(d[15]), .s(n17687), .op(n13545) );
  mux2_1 U21477 ( .ip1(\LUT[4][14] ), .ip2(d[14]), .s(n17687), .op(n13544) );
  mux2_1 U21478 ( .ip1(\LUT[4][13] ), .ip2(d[13]), .s(n17687), .op(n13543) );
  mux2_1 U21479 ( .ip1(\LUT[4][12] ), .ip2(d[12]), .s(n17687), .op(n13542) );
  mux2_1 U21480 ( .ip1(\LUT[4][11] ), .ip2(d[11]), .s(n17687), .op(n13541) );
  mux2_1 U21481 ( .ip1(\LUT[4][10] ), .ip2(d[10]), .s(n17687), .op(n13540) );
  mux2_1 U21482 ( .ip1(\LUT[4][9] ), .ip2(d[9]), .s(n17687), .op(n13539) );
  mux2_1 U21483 ( .ip1(\LUT[4][8] ), .ip2(d[8]), .s(n17687), .op(n13538) );
  mux2_1 U21484 ( .ip1(\LUT[4][7] ), .ip2(d[7]), .s(n17687), .op(n13537) );
  mux2_1 U21485 ( .ip1(\LUT[4][6] ), .ip2(d[6]), .s(n17687), .op(n13536) );
  mux2_1 U21486 ( .ip1(\LUT[4][5] ), .ip2(d[5]), .s(n17688), .op(n13535) );
  mux2_1 U21487 ( .ip1(\LUT[4][4] ), .ip2(d[4]), .s(n17688), .op(n13534) );
  mux2_1 U21488 ( .ip1(\LUT[4][3] ), .ip2(d[3]), .s(n17688), .op(n13533) );
  mux2_1 U21489 ( .ip1(\LUT[4][2] ), .ip2(d[2]), .s(n17688), .op(n13532) );
  mux2_1 U21490 ( .ip1(\LUT[4][1] ), .ip2(d[1]), .s(n17688), .op(n13531) );
  mux2_1 U21491 ( .ip1(\LUT[4][0] ), .ip2(d[0]), .s(n17688), .op(n13530) );
  mux2_1 U21492 ( .ip1(\LUT[3][15] ), .ip2(n17629), .s(n17689), .op(n13529) );
  mux2_1 U21493 ( .ip1(\LUT[3][14] ), .ip2(n17630), .s(n17689), .op(n13528) );
  mux2_1 U21494 ( .ip1(\LUT[3][13] ), .ip2(n17631), .s(n17689), .op(n13527) );
  mux2_1 U21495 ( .ip1(\LUT[3][12] ), .ip2(n17632), .s(n17689), .op(n13526) );
  mux2_1 U21496 ( .ip1(\LUT[3][11] ), .ip2(n17633), .s(n17689), .op(n13525) );
  mux2_1 U21497 ( .ip1(\LUT[3][10] ), .ip2(n17634), .s(n17689), .op(n13524) );
  mux2_1 U21498 ( .ip1(\LUT[3][9] ), .ip2(n17635), .s(n17689), .op(n13523) );
  mux2_1 U21499 ( .ip1(\LUT[3][8] ), .ip2(n17636), .s(n17689), .op(n13522) );
  mux2_1 U21500 ( .ip1(\LUT[3][7] ), .ip2(n17637), .s(n17689), .op(n13521) );
  mux2_1 U21501 ( .ip1(\LUT[3][6] ), .ip2(n17639), .s(n17689), .op(n13520) );
  mux2_1 U21502 ( .ip1(\LUT[3][5] ), .ip2(n17640), .s(n17690), .op(n13519) );
  mux2_1 U21503 ( .ip1(\LUT[3][4] ), .ip2(n17641), .s(n17690), .op(n13518) );
  mux2_1 U21504 ( .ip1(\LUT[3][3] ), .ip2(n17642), .s(n17690), .op(n13517) );
  mux2_1 U21505 ( .ip1(\LUT[3][2] ), .ip2(n17643), .s(n17690), .op(n13516) );
  mux2_1 U21506 ( .ip1(\LUT[3][1] ), .ip2(n17644), .s(n17690), .op(n13515) );
  mux2_1 U21507 ( .ip1(\LUT[3][0] ), .ip2(n17646), .s(n17690), .op(n13514) );
  mux2_1 U21508 ( .ip1(\LUT[2][15] ), .ip2(d[15]), .s(n17691), .op(n13513) );
  mux2_1 U21509 ( .ip1(\LUT[2][14] ), .ip2(d[14]), .s(n17691), .op(n13512) );
  mux2_1 U21510 ( .ip1(\LUT[2][13] ), .ip2(d[13]), .s(n17691), .op(n13511) );
  mux2_1 U21511 ( .ip1(\LUT[2][12] ), .ip2(d[12]), .s(n17691), .op(n13510) );
  mux2_1 U21512 ( .ip1(\LUT[2][11] ), .ip2(d[11]), .s(n17691), .op(n13509) );
  mux2_1 U21513 ( .ip1(\LUT[2][10] ), .ip2(d[10]), .s(n17691), .op(n13508) );
  mux2_1 U21514 ( .ip1(\LUT[2][9] ), .ip2(d[9]), .s(n17691), .op(n13507) );
  mux2_1 U21515 ( .ip1(\LUT[2][8] ), .ip2(d[8]), .s(n17691), .op(n13506) );
  mux2_1 U21516 ( .ip1(\LUT[2][7] ), .ip2(d[7]), .s(n17691), .op(n13505) );
  mux2_1 U21517 ( .ip1(\LUT[2][6] ), .ip2(d[6]), .s(n17691), .op(n13504) );
  mux2_1 U21518 ( .ip1(\LUT[2][5] ), .ip2(d[5]), .s(n17692), .op(n13503) );
  mux2_1 U21519 ( .ip1(\LUT[2][4] ), .ip2(d[4]), .s(n17692), .op(n13502) );
  mux2_1 U21520 ( .ip1(\LUT[2][3] ), .ip2(d[3]), .s(n17692), .op(n13501) );
  mux2_1 U21521 ( .ip1(\LUT[2][2] ), .ip2(d[2]), .s(n17692), .op(n13500) );
  mux2_1 U21522 ( .ip1(\LUT[2][1] ), .ip2(d[1]), .s(n17692), .op(n13499) );
  mux2_1 U21523 ( .ip1(\LUT[2][0] ), .ip2(d[0]), .s(n17692), .op(n13498) );
  mux2_1 U21524 ( .ip1(\LUT[1][15] ), .ip2(d[15]), .s(n17693), .op(n13497) );
  mux2_1 U21525 ( .ip1(\LUT[1][14] ), .ip2(d[14]), .s(n17693), .op(n13496) );
  mux2_1 U21526 ( .ip1(\LUT[1][13] ), .ip2(d[13]), .s(n17693), .op(n13495) );
  mux2_1 U21527 ( .ip1(\LUT[1][12] ), .ip2(d[12]), .s(n17693), .op(n13494) );
  mux2_1 U21528 ( .ip1(\LUT[1][11] ), .ip2(d[11]), .s(n17693), .op(n13493) );
  mux2_1 U21529 ( .ip1(\LUT[1][10] ), .ip2(d[10]), .s(n17693), .op(n13492) );
  mux2_1 U21530 ( .ip1(\LUT[1][9] ), .ip2(d[9]), .s(n17693), .op(n13491) );
  mux2_1 U21531 ( .ip1(\LUT[1][8] ), .ip2(d[8]), .s(n17693), .op(n13490) );
  mux2_1 U21532 ( .ip1(\LUT[1][7] ), .ip2(d[7]), .s(n17693), .op(n13489) );
  mux2_1 U21533 ( .ip1(\LUT[1][6] ), .ip2(d[6]), .s(n17693), .op(n13488) );
  mux2_1 U21534 ( .ip1(\LUT[1][5] ), .ip2(d[5]), .s(n17694), .op(n13487) );
  mux2_1 U21535 ( .ip1(\LUT[1][4] ), .ip2(d[4]), .s(n17694), .op(n13486) );
  mux2_1 U21536 ( .ip1(\LUT[1][3] ), .ip2(d[3]), .s(n17694), .op(n13485) );
  mux2_1 U21537 ( .ip1(\LUT[1][2] ), .ip2(d[2]), .s(n17694), .op(n13484) );
  mux2_1 U21538 ( .ip1(\LUT[1][1] ), .ip2(d[1]), .s(n17694), .op(n13483) );
  mux2_1 U21539 ( .ip1(\LUT[1][0] ), .ip2(d[0]), .s(n17694), .op(n13482) );
  mux2_1 U21540 ( .ip1(\LUT[0][15] ), .ip2(d[15]), .s(n17695), .op(n13481) );
  mux2_1 U21541 ( .ip1(\LUT[0][14] ), .ip2(d[14]), .s(n17695), .op(n13480) );
  mux2_1 U21542 ( .ip1(\LUT[0][13] ), .ip2(d[13]), .s(n17695), .op(n13479) );
  mux2_1 U21543 ( .ip1(\LUT[0][12] ), .ip2(d[12]), .s(n17695), .op(n13478) );
  mux2_1 U21544 ( .ip1(\LUT[0][11] ), .ip2(d[11]), .s(n17695), .op(n13477) );
  mux2_1 U21545 ( .ip1(\LUT[0][10] ), .ip2(d[10]), .s(n17695), .op(n13476) );
  mux2_1 U21546 ( .ip1(\LUT[0][9] ), .ip2(d[9]), .s(n17695), .op(n13475) );
  mux2_1 U21547 ( .ip1(\LUT[0][8] ), .ip2(d[8]), .s(n17695), .op(n13474) );
  mux2_1 U21548 ( .ip1(\LUT[0][7] ), .ip2(d[7]), .s(n17695), .op(n13473) );
  mux2_1 U21549 ( .ip1(\LUT[0][6] ), .ip2(d[6]), .s(n17695), .op(n13472) );
  mux2_1 U21550 ( .ip1(\LUT[0][5] ), .ip2(d[5]), .s(n17696), .op(n13471) );
  mux2_1 U21551 ( .ip1(\LUT[0][4] ), .ip2(d[4]), .s(n17696), .op(n13470) );
  mux2_1 U21552 ( .ip1(\LUT[0][3] ), .ip2(d[3]), .s(n17696), .op(n13469) );
  mux2_1 U21553 ( .ip1(\LUT[0][2] ), .ip2(d[2]), .s(n17696), .op(n13468) );
  mux2_1 U21554 ( .ip1(\LUT[0][1] ), .ip2(d[1]), .s(n17696), .op(n13467) );
  mux2_1 U21555 ( .ip1(\LUT[0][0] ), .ip2(d[0]), .s(n17696), .op(n13466) );
  nor4_1 U21556 ( .ip1(sig_in[14]), .ip2(n17981), .ip3(n17845), .ip4(
        sig_in[13]), .op(n17697) );
  or2_1 U21557 ( .ip1(n17697), .ip2(sig_in[15]), .op(n17703) );
  inv_1 U21558 ( .ip(n20652), .op(n24464) );
  nor3_1 U21559 ( .ip1(sig_in[2]), .ip2(n24464), .ip3(sig_in[8]), .op(n17699)
         );
  buf_1 U21560 ( .ip(sig_in[7]), .op(n17732) );
  nor4_1 U21561 ( .ip1(sig_in[0]), .ip2(sig_in[3]), .ip3(sig_in[6]), .ip4(
        n17732), .op(n17698) );
  buf_1 U21562 ( .ip(sig_in[4]), .op(n24462) );
  buf_1 U21563 ( .ip(sig_in[5]), .op(n22833) );
  nand4_1 U21564 ( .ip1(n17699), .ip2(n17698), .ip3(n23721), .ip4(n23283), 
        .op(n17700) );
  nand3_1 U21565 ( .ip1(sig_in[10]), .ip2(sig_in[9]), .ip3(n17700), .op(n17701) );
  or2_1 U21566 ( .ip1(n17701), .ip2(sig_in[15]), .op(n17702) );
  nand2_1 U21567 ( .ip1(n17703), .ip2(n17702), .op(n26294) );
  or2_1 U21568 ( .ip1(sig_in[15]), .ip2(n26294), .op(n17707) );
  inv_1 U21569 ( .ip(sig_in[10]), .op(n24370) );
  inv_1 U21570 ( .ip(n17845), .op(n24233) );
  inv_1 U21571 ( .ip(sig_in[13]), .op(n24332) );
  not_ab_or_c_or_d U21572 ( .ip1(n24269), .ip2(n23980), .ip3(n24233), .ip4(
        n24376), .op(n17704) );
  nand3_1 U21573 ( .ip1(sig_in[14]), .ip2(n17981), .ip3(n17704), .op(n17705)
         );
  or2_1 U21574 ( .ip1(n17705), .ip2(n26294), .op(n17706) );
  nand2_1 U21575 ( .ip1(n17707), .ip2(n17706), .op(n24518) );
  inv_1 U21576 ( .ip(n24518), .op(n24521) );
  inv_1 U21577 ( .ip(sig_in[15]), .op(n24329) );
  buf_1 U21578 ( .ip(n24329), .op(n24090) );
  nor2_1 U21579 ( .ip1(\x[29][15] ), .ip2(n24090), .op(n17760) );
  nor3_1 U21580 ( .ip1(n17760), .ip2(\x[29][14] ), .ip3(n24382), .op(n17708)
         );
  or2_1 U21581 ( .ip1(\x[29][15] ), .ip2(n17708), .op(n17710) );
  or2_1 U21582 ( .ip1(n24180), .ip2(n17708), .op(n17709) );
  nand2_1 U21583 ( .ip1(n17710), .ip2(n17709), .op(n24222) );
  inv_1 U21584 ( .ip(sig_in[14]), .op(n24230) );
  buf_1 U21585 ( .ip(n24230), .op(n24327) );
  nor2_1 U21586 ( .ip1(\x[30][14] ), .ip2(n24327), .op(n17711) );
  or2_1 U21587 ( .ip1(\x[30][15] ), .ip2(n17711), .op(n17713) );
  or2_1 U21588 ( .ip1(n24180), .ip2(n17711), .op(n17712) );
  nand2_1 U21589 ( .ip1(n17713), .ip2(n17712), .op(n17759) );
  buf_1 U21590 ( .ip(n24332), .op(n24235) );
  buf_1 U21591 ( .ip(n24235), .op(n24081) );
  nand2_1 U21592 ( .ip1(\x[30][13] ), .ip2(n24081), .op(n17715) );
  nand2_1 U21593 ( .ip1(\x[30][14] ), .ip2(n24327), .op(n17714) );
  nand2_1 U21594 ( .ip1(n17715), .ip2(n17714), .op(n17758) );
  nor2_1 U21595 ( .ip1(\x[30][15] ), .ip2(n24090), .op(n17757) );
  inv_1 U21596 ( .ip(n17981), .op(n24136) );
  not_ab_or_c_or_d U21597 ( .ip1(\x[30][11] ), .ip2(n24136), .ip3(\x[30][10] ), 
        .ip4(n23980), .op(n17749) );
  nor2_1 U21598 ( .ip1(\x[30][7] ), .ip2(n24142), .op(n17738) );
  inv_1 U21599 ( .ip(sig_in[8]), .op(n24358) );
  nor2_1 U21600 ( .ip1(\x[30][8] ), .ip2(n24358), .op(n17737) );
  inv_1 U21601 ( .ip(n24455), .op(n21171) );
  inv_1 U21602 ( .ip(n21171), .op(n24043) );
  nor2_1 U21603 ( .ip1(\x[30][9] ), .ip2(n24043), .op(n17739) );
  inv_1 U21604 ( .ip(sig_in[5]), .op(n23600) );
  and2_1 U21605 ( .ip1(n24045), .ip2(\x[30][6] ), .op(n17729) );
  inv_1 U21606 ( .ip(\x[30][4] ), .op(n17727) );
  nor2_1 U21607 ( .ip1(n24462), .ip2(n17727), .op(n17724) );
  inv_1 U21608 ( .ip(\x[30][3] ), .op(n17722) );
  inv_1 U21609 ( .ip(sig_in[2]), .op(n24107) );
  inv_1 U21610 ( .ip(n20652), .op(n22513) );
  inv_1 U21611 ( .ip(\x[30][1] ), .op(n17717) );
  nor2_1 U21612 ( .ip1(n22513), .ip2(n17717), .op(n17719) );
  inv_1 U21613 ( .ip(n20652), .op(n24467) );
  inv_1 U21614 ( .ip(\x[30][0] ), .op(n17716) );
  not_ab_or_c_or_d U21615 ( .ip1(n24467), .ip2(n17717), .ip3(sig_in[0]), .ip4(
        n17716), .op(n17718) );
  not_ab_or_c_or_d U21616 ( .ip1(\x[30][2] ), .ip2(n24335), .ip3(n17719), 
        .ip4(n17718), .op(n17721) );
  buf_1 U21617 ( .ip(n24107), .op(n24463) );
  nor2_1 U21618 ( .ip1(\x[30][2] ), .ip2(n24463), .op(n17720) );
  not_ab_or_c_or_d U21619 ( .ip1(sig_in[3]), .ip2(n17722), .ip3(n17721), .ip4(
        n17720), .op(n17723) );
  not_ab_or_c_or_d U21620 ( .ip1(\x[30][3] ), .ip2(n22795), .ip3(n17724), 
        .ip4(n17723), .op(n17726) );
  inv_1 U21621 ( .ip(n22833), .op(n23283) );
  buf_1 U21622 ( .ip(n23283), .op(n24350) );
  nor2_1 U21623 ( .ip1(\x[30][5] ), .ip2(n24350), .op(n17725) );
  not_ab_or_c_or_d U21624 ( .ip1(sig_in[4]), .ip2(n17727), .ip3(n17726), .ip4(
        n17725), .op(n17728) );
  not_ab_or_c_or_d U21625 ( .ip1(\x[30][5] ), .ip2(n23600), .ip3(n17729), 
        .ip4(n17728), .op(n17731) );
  inv_1 U21626 ( .ip(sig_in[6]), .op(n23509) );
  nor2_1 U21627 ( .ip1(\x[30][6] ), .ip2(n23509), .op(n17730) );
  nor2_1 U21628 ( .ip1(n17731), .ip2(n17730), .op(n17733) );
  or2_1 U21629 ( .ip1(\x[30][7] ), .ip2(n17733), .op(n17735) );
  or2_1 U21630 ( .ip1(n24044), .ip2(n17733), .op(n17734) );
  nand2_1 U21631 ( .ip1(n17735), .ip2(n17734), .op(n17736) );
  nor4_1 U21632 ( .ip1(n17738), .ip2(n17737), .ip3(n17739), .ip4(n17736), .op(
        n17745) );
  nand2_1 U21633 ( .ip1(\x[30][11] ), .ip2(n21793), .op(n17743) );
  inv_1 U21634 ( .ip(n17739), .op(n17740) );
  nand3_1 U21635 ( .ip1(\x[30][8] ), .ip2(n23804), .ip3(n17740), .op(n17742)
         );
  buf_1 U21636 ( .ip(n24370), .op(n23980) );
  nand2_1 U21637 ( .ip1(\x[30][10] ), .ip2(n23980), .op(n17741) );
  nand3_1 U21638 ( .ip1(n17743), .ip2(n17742), .ip3(n17741), .op(n17744) );
  not_ab_or_c_or_d U21639 ( .ip1(\x[30][9] ), .ip2(n24269), .ip3(n17745), 
        .ip4(n17744), .op(n17748) );
  inv_1 U21640 ( .ip(n17845), .op(n24449) );
  nor2_1 U21641 ( .ip1(\x[30][12] ), .ip2(n24449), .op(n17747) );
  nor2_1 U21642 ( .ip1(\x[30][11] ), .ip2(n21793), .op(n17746) );
  or4_1 U21643 ( .ip1(n17749), .ip2(n17748), .ip3(n17747), .ip4(n17746), .op(
        n17751) );
  or2_1 U21644 ( .ip1(n24137), .ip2(\x[30][13] ), .op(n17750) );
  nand2_1 U21645 ( .ip1(n17759), .ip2(n17750), .op(n17752) );
  or2_1 U21646 ( .ip1(n17751), .ip2(n17752), .op(n17755) );
  buf_1 U21647 ( .ip(sig_in[12]), .op(n17845) );
  nand2_1 U21648 ( .ip1(\x[30][12] ), .ip2(n24079), .op(n17753) );
  or2_1 U21649 ( .ip1(n17753), .ip2(n17752), .op(n17754) );
  nand2_1 U21650 ( .ip1(n17755), .ip2(n17754), .op(n17756) );
  not_ab_or_c_or_d U21651 ( .ip1(n17759), .ip2(n17758), .ip3(n17757), .ip4(
        n17756), .op(n18494) );
  or2_1 U21652 ( .ip1(n24222), .ip2(n18494), .op(n17809) );
  buf_1 U21653 ( .ip(n24230), .op(n23938) );
  nand2_1 U21654 ( .ip1(n23938), .ip2(\x[29][14] ), .op(n17763) );
  inv_1 U21655 ( .ip(n17760), .op(n17762) );
  nand2_1 U21656 ( .ip1(\x[29][13] ), .ip2(n24081), .op(n17761) );
  nand3_1 U21657 ( .ip1(n17763), .ip2(n17762), .ip3(n17761), .op(n24218) );
  or2_1 U21658 ( .ip1(\x[29][12] ), .ip2(n24218), .op(n17765) );
  or2_1 U21659 ( .ip1(n24449), .ip2(n24218), .op(n17764) );
  nand2_1 U21660 ( .ip1(n17765), .ip2(n17764), .op(n24226) );
  nor2_1 U21661 ( .ip1(\x[29][13] ), .ip2(n23895), .op(n17766) );
  or2_1 U21662 ( .ip1(sig_in[12]), .ip2(n17766), .op(n17769) );
  inv_1 U21663 ( .ip(\x[29][12] ), .op(n17767) );
  or2_1 U21664 ( .ip1(n17767), .ip2(n17766), .op(n17768) );
  nand2_1 U21665 ( .ip1(n17769), .ip2(n17768), .op(n24217) );
  inv_1 U21666 ( .ip(\x[29][11] ), .op(n17805) );
  buf_1 U21667 ( .ip(n24370), .op(n20880) );
  nor2_1 U21668 ( .ip1(\x[29][10] ), .ip2(n20880), .op(n17770) );
  or2_1 U21669 ( .ip1(sig_in[9]), .ip2(n17770), .op(n17773) );
  inv_1 U21670 ( .ip(\x[29][9] ), .op(n17771) );
  or2_1 U21671 ( .ip1(n17771), .ip2(n17770), .op(n17772) );
  nand2_1 U21672 ( .ip1(n17773), .ip2(n17772), .op(n17776) );
  nand2_1 U21673 ( .ip1(\x[29][10] ), .ip2(n23980), .op(n17775) );
  inv_1 U21674 ( .ip(n17981), .op(n24456) );
  nand2_1 U21675 ( .ip1(\x[29][11] ), .ip2(n24456), .op(n17774) );
  nand2_1 U21676 ( .ip1(n17775), .ip2(n17774), .op(n17796) );
  nor2_1 U21677 ( .ip1(n17776), .ip2(n17796), .op(n17804) );
  inv_1 U21678 ( .ip(n17732), .op(n24461) );
  and2_1 U21679 ( .ip1(n24461), .ip2(\x[29][7] ), .op(n17793) );
  inv_1 U21680 ( .ip(\x[29][5] ), .op(n17791) );
  nor2_1 U21681 ( .ip1(sig_in[5]), .ip2(n17791), .op(n17788) );
  inv_1 U21682 ( .ip(n24462), .op(n23721) );
  nor2_1 U21683 ( .ip1(\x[29][4] ), .ip2(n23721), .op(n17786) );
  inv_1 U21684 ( .ip(sig_in[3]), .op(n24342) );
  buf_1 U21685 ( .ip(n24107), .op(n24470) );
  not_ab_or_c_or_d U21686 ( .ip1(\x[29][3] ), .ip2(n24342), .ip3(\x[29][2] ), 
        .ip4(n24470), .op(n17785) );
  nor2_1 U21687 ( .ip1(\x[29][3] ), .ip2(n22525), .op(n17784) );
  inv_1 U21688 ( .ip(\x[29][1] ), .op(n17778) );
  inv_1 U21689 ( .ip(\x[29][0] ), .op(n17777) );
  not_ab_or_c_or_d U21690 ( .ip1(n22513), .ip2(n17778), .ip3(sig_in[0]), .ip4(
        n17777), .op(n17782) );
  nand2_1 U21691 ( .ip1(\x[29][3] ), .ip2(n22795), .op(n17780) );
  nand2_1 U21692 ( .ip1(\x[29][1] ), .ip2(n21685), .op(n17779) );
  nand2_1 U21693 ( .ip1(n17780), .ip2(n17779), .op(n17781) );
  not_ab_or_c_or_d U21694 ( .ip1(\x[29][2] ), .ip2(n24470), .ip3(n17782), 
        .ip4(n17781), .op(n17783) );
  nor4_1 U21695 ( .ip1(n17786), .ip2(n17785), .ip3(n17784), .ip4(n17783), .op(
        n17787) );
  not_ab_or_c_or_d U21696 ( .ip1(\x[29][4] ), .ip2(n24256), .ip3(n17788), 
        .ip4(n17787), .op(n17790) );
  inv_1 U21697 ( .ip(sig_in[6]), .op(n24485) );
  nor2_1 U21698 ( .ip1(\x[29][6] ), .ip2(n24485), .op(n17789) );
  not_ab_or_c_or_d U21699 ( .ip1(n22833), .ip2(n17791), .ip3(n17790), .ip4(
        n17789), .op(n17792) );
  not_ab_or_c_or_d U21700 ( .ip1(\x[29][6] ), .ip2(n24485), .ip3(n17793), 
        .ip4(n17792), .op(n17795) );
  inv_1 U21701 ( .ip(n17732), .op(n24492) );
  nor2_1 U21702 ( .ip1(\x[29][7] ), .ip2(n24492), .op(n17794) );
  nor2_1 U21703 ( .ip1(n17795), .ip2(n17794), .op(n17800) );
  inv_1 U21704 ( .ip(n17796), .op(n17798) );
  nand2_1 U21705 ( .ip1(\x[29][9] ), .ip2(n24269), .op(n17797) );
  nand2_1 U21706 ( .ip1(n17798), .ip2(n17797), .op(n17799) );
  nor3_1 U21707 ( .ip1(n17800), .ip2(\x[29][8] ), .ip3(n17799), .op(n17802) );
  inv_1 U21708 ( .ip(sig_in[8]), .op(n24491) );
  not_ab_or_c_or_d U21709 ( .ip1(n17800), .ip2(\x[29][8] ), .ip3(n24491), 
        .ip4(n17799), .op(n17801) );
  or2_1 U21710 ( .ip1(n17802), .ip2(n17801), .op(n17803) );
  not_ab_or_c_or_d U21711 ( .ip1(sig_in[11]), .ip2(n17805), .ip3(n17804), 
        .ip4(n17803), .op(n24194) );
  nand2_1 U21712 ( .ip1(n24217), .ip2(n24194), .op(n17806) );
  nand2_1 U21713 ( .ip1(n24226), .ip2(n17806), .op(n17807) );
  or2_1 U21714 ( .ip1(n17807), .ip2(n18494), .op(n17808) );
  nand2_1 U21715 ( .ip1(n17809), .ip2(n17808), .op(n24850) );
  buf_1 U21716 ( .ip(n24329), .op(n24186) );
  nand2_1 U21717 ( .ip1(\x[34][15] ), .ip2(n24186), .op(n18439) );
  inv_1 U21718 ( .ip(sig_in[14]), .op(n24185) );
  or2_1 U21719 ( .ip1(n24185), .ip2(\x[34][14] ), .op(n17810) );
  nand2_1 U21720 ( .ip1(n18439), .ip2(n17810), .op(n18447) );
  or2_1 U21721 ( .ip1(n24180), .ip2(\x[34][15] ), .op(n17893) );
  inv_1 U21722 ( .ip(n17845), .op(n24079) );
  nor2_1 U21723 ( .ip1(\x[34][12] ), .ip2(n24079), .op(n17844) );
  nor2_1 U21724 ( .ip1(\x[34][11] ), .ip2(n24456), .op(n17843) );
  nor2_1 U21725 ( .ip1(\x[34][13] ), .ip2(n24332), .op(n17842) );
  inv_1 U21726 ( .ip(n17981), .op(n24371) );
  and2_1 U21727 ( .ip1(n24371), .ip2(\x[34][11] ), .op(n17838) );
  nor3_1 U21728 ( .ip1(n20880), .ip2(\x[34][10] ), .ip3(n17838), .op(n17840)
         );
  inv_1 U21729 ( .ip(sig_in[9]), .op(n24455) );
  nor2_1 U21730 ( .ip1(\x[34][9] ), .ip2(n24455), .op(n17836) );
  and2_1 U21731 ( .ip1(n24100), .ip2(\x[34][8] ), .op(n17834) );
  inv_1 U21732 ( .ip(\x[34][7] ), .op(n17831) );
  nor2_1 U21733 ( .ip1(\x[34][8] ), .ip2(n24358), .op(n17830) );
  inv_1 U21734 ( .ip(sig_in[6]), .op(n24045) );
  nor2_1 U21735 ( .ip1(n17732), .ip2(n17831), .op(n17826) );
  nor3_1 U21736 ( .ip1(n24045), .ip2(\x[34][6] ), .ip3(n17826), .op(n17828) );
  nor2_1 U21737 ( .ip1(\x[34][5] ), .ip2(n23283), .op(n17824) );
  and2_1 U21738 ( .ip1(n23860), .ip2(\x[34][4] ), .op(n17822) );
  inv_1 U21739 ( .ip(\x[34][3] ), .op(n17819) );
  buf_1 U21740 ( .ip(n24107), .op(n24335) );
  and2_1 U21741 ( .ip1(n24335), .ip2(\x[34][2] ), .op(n17816) );
  nand2_1 U21742 ( .ip1(\x[34][1] ), .ip2(n20652), .op(n17814) );
  nand2_1 U21743 ( .ip1(\x[34][0] ), .ip2(n24143), .op(n17813) );
  nor2_1 U21744 ( .ip1(\x[34][2] ), .ip2(n24463), .op(n17812) );
  nor2_1 U21745 ( .ip1(\x[34][1] ), .ip2(n21685), .op(n17811) );
  not_ab_or_c_or_d U21746 ( .ip1(n17814), .ip2(n17813), .ip3(n17812), .ip4(
        n17811), .op(n17815) );
  not_ab_or_c_or_d U21747 ( .ip1(\x[34][3] ), .ip2(n22795), .ip3(n17816), 
        .ip4(n17815), .op(n17818) );
  inv_1 U21748 ( .ip(n24462), .op(n24256) );
  nor2_1 U21749 ( .ip1(\x[34][4] ), .ip2(n24256), .op(n17817) );
  not_ab_or_c_or_d U21750 ( .ip1(n23251), .ip2(n17819), .ip3(n17818), .ip4(
        n17817), .op(n17821) );
  and2_1 U21751 ( .ip1(n23283), .ip2(\x[34][5] ), .op(n17820) );
  nor3_1 U21752 ( .ip1(n17822), .ip2(n17821), .ip3(n17820), .op(n17823) );
  nor2_1 U21753 ( .ip1(n17824), .ip2(n17823), .op(n17825) );
  not_ab_or_c_or_d U21754 ( .ip1(\x[34][6] ), .ip2(n23509), .ip3(n17826), 
        .ip4(n17825), .op(n17827) );
  or2_1 U21755 ( .ip1(n17828), .ip2(n17827), .op(n17829) );
  not_ab_or_c_or_d U21756 ( .ip1(sig_in[7]), .ip2(n17831), .ip3(n17830), .ip4(
        n17829), .op(n17833) );
  and2_1 U21757 ( .ip1(n24269), .ip2(\x[34][9] ), .op(n17832) );
  nor3_1 U21758 ( .ip1(n17834), .ip2(n17833), .ip3(n17832), .op(n17835) );
  nor2_1 U21759 ( .ip1(n17836), .ip2(n17835), .op(n17837) );
  not_ab_or_c_or_d U21760 ( .ip1(\x[34][10] ), .ip2(n23980), .ip3(n17838), 
        .ip4(n17837), .op(n17839) );
  or2_1 U21761 ( .ip1(n17840), .ip2(n17839), .op(n17841) );
  nor4_1 U21762 ( .ip1(n17844), .ip2(n17843), .ip3(n17842), .ip4(n17841), .op(
        n18444) );
  nand2_1 U21763 ( .ip1(\x[34][13] ), .ip2(n24235), .op(n17847) );
  nand2_1 U21764 ( .ip1(\x[34][12] ), .ip2(n24233), .op(n17846) );
  nand2_1 U21765 ( .ip1(n17847), .ip2(n17846), .op(n18445) );
  nand2_1 U21766 ( .ip1(\x[34][14] ), .ip2(n24230), .op(n17848) );
  nand2_1 U21767 ( .ip1(n17893), .ip2(n17848), .op(n18438) );
  nor3_1 U21768 ( .ip1(n18444), .ip2(n18445), .ip3(n18438), .op(n17892) );
  buf_1 U21769 ( .ip(n24329), .op(n24384) );
  nor2_1 U21770 ( .ip1(n24384), .ip2(\x[33][15] ), .op(n17890) );
  buf_1 U21771 ( .ip(n24332), .op(n23895) );
  and2_1 U21772 ( .ip1(n23895), .ip2(\x[33][13] ), .op(n17881) );
  and2_1 U21773 ( .ip1(n24461), .ip2(\x[33][7] ), .op(n17865) );
  inv_1 U21774 ( .ip(\x[33][3] ), .op(n17855) );
  nor2_1 U21775 ( .ip1(\x[33][2] ), .ip2(n24463), .op(n17854) );
  inv_1 U21776 ( .ip(\x[33][1] ), .op(n17850) );
  nor2_1 U21777 ( .ip1(n22513), .ip2(n17850), .op(n17852) );
  inv_1 U21778 ( .ip(\x[33][0] ), .op(n17849) );
  not_ab_or_c_or_d U21779 ( .ip1(n24464), .ip2(n17850), .ip3(sig_in[0]), .ip4(
        n17849), .op(n17851) );
  not_ab_or_c_or_d U21780 ( .ip1(\x[33][2] ), .ip2(n24335), .ip3(n17852), 
        .ip4(n17851), .op(n17853) );
  not_ab_or_c_or_d U21781 ( .ip1(n23251), .ip2(n17855), .ip3(n17854), .ip4(
        n17853), .op(n17859) );
  nand2_1 U21782 ( .ip1(\x[33][5] ), .ip2(n23283), .op(n17857) );
  nand2_1 U21783 ( .ip1(\x[33][4] ), .ip2(n23860), .op(n17856) );
  nand2_1 U21784 ( .ip1(n17857), .ip2(n17856), .op(n17858) );
  not_ab_or_c_or_d U21785 ( .ip1(\x[33][3] ), .ip2(n22795), .ip3(n17859), 
        .ip4(n17858), .op(n17863) );
  nor2_1 U21786 ( .ip1(\x[33][5] ), .ip2(n23283), .op(n17862) );
  nor2_1 U21787 ( .ip1(\x[33][6] ), .ip2(n24485), .op(n17861) );
  buf_1 U21788 ( .ip(n23600), .op(n24482) );
  inv_1 U21789 ( .ip(n24462), .op(n24347) );
  not_ab_or_c_or_d U21790 ( .ip1(\x[33][5] ), .ip2(n24482), .ip3(\x[33][4] ), 
        .ip4(n24347), .op(n17860) );
  nor4_1 U21791 ( .ip1(n17863), .ip2(n17862), .ip3(n17861), .ip4(n17860), .op(
        n17864) );
  not_ab_or_c_or_d U21792 ( .ip1(\x[33][6] ), .ip2(n23509), .ip3(n17865), 
        .ip4(n17864), .op(n17868) );
  nor2_1 U21793 ( .ip1(\x[33][9] ), .ip2(n24043), .op(n17869) );
  inv_1 U21794 ( .ip(sig_in[8]), .op(n23971) );
  nor2_1 U21795 ( .ip1(\x[33][8] ), .ip2(n23971), .op(n17867) );
  inv_1 U21796 ( .ip(n17732), .op(n24142) );
  nor2_1 U21797 ( .ip1(\x[33][7] ), .ip2(n24142), .op(n17866) );
  nor4_1 U21798 ( .ip1(n17868), .ip2(n17869), .ip3(n17867), .ip4(n17866), .op(
        n17875) );
  nand2_1 U21799 ( .ip1(n24370), .ip2(\x[33][10] ), .op(n17873) );
  inv_1 U21800 ( .ip(n17869), .op(n17870) );
  nand3_1 U21801 ( .ip1(\x[33][8] ), .ip2(n24100), .ip3(n17870), .op(n17872)
         );
  nand2_1 U21802 ( .ip1(\x[33][11] ), .ip2(n21793), .op(n17871) );
  nand3_1 U21803 ( .ip1(n17873), .ip2(n17872), .ip3(n17871), .op(n17874) );
  not_ab_or_c_or_d U21804 ( .ip1(\x[33][9] ), .ip2(n24164), .ip3(n17875), 
        .ip4(n17874), .op(n17879) );
  nor2_1 U21805 ( .ip1(\x[33][11] ), .ip2(n21793), .op(n17878) );
  nor2_1 U21806 ( .ip1(\x[33][12] ), .ip2(n24079), .op(n17877) );
  not_ab_or_c_or_d U21807 ( .ip1(\x[33][11] ), .ip2(n24136), .ip3(\x[33][10] ), 
        .ip4(n23980), .op(n17876) );
  nor4_1 U21808 ( .ip1(n17879), .ip2(n17878), .ip3(n17877), .ip4(n17876), .op(
        n17880) );
  not_ab_or_c_or_d U21809 ( .ip1(\x[33][12] ), .ip2(n24079), .ip3(n17881), 
        .ip4(n17880), .op(n17883) );
  nor2_1 U21810 ( .ip1(\x[33][13] ), .ip2(n24332), .op(n17882) );
  nor2_1 U21811 ( .ip1(n17883), .ip2(n17882), .op(n17884) );
  or2_1 U21812 ( .ip1(\x[33][14] ), .ip2(n17884), .op(n17886) );
  buf_1 U21813 ( .ip(n24185), .op(n24382) );
  or2_1 U21814 ( .ip1(n24382), .ip2(n17884), .op(n17885) );
  nand2_1 U21815 ( .ip1(n17886), .ip2(n17885), .op(n17888) );
  nor2_1 U21816 ( .ip1(\x[33][14] ), .ip2(n24327), .op(n17887) );
  not_ab_or_c_or_d U21817 ( .ip1(\x[33][15] ), .ip2(n24180), .ip3(n17888), 
        .ip4(n17887), .op(n17889) );
  nor2_1 U21818 ( .ip1(n17890), .ip2(n17889), .op(n17937) );
  inv_1 U21819 ( .ip(n17937), .op(n17891) );
  not_ab_or_c_or_d U21820 ( .ip1(n18447), .ip2(n17893), .ip3(n17892), .ip4(
        n17891), .op(n24889) );
  nand2_1 U21821 ( .ip1(\x[32][15] ), .ip2(n24186), .op(n17938) );
  or2_1 U21822 ( .ip1(n24180), .ip2(\x[32][15] ), .op(n18504) );
  nand2_1 U21823 ( .ip1(\x[32][14] ), .ip2(n23938), .op(n17894) );
  nand2_1 U21824 ( .ip1(n18504), .ip2(n17894), .op(n18498) );
  and2_1 U21825 ( .ip1(n23895), .ip2(\x[32][13] ), .op(n17895) );
  or2_1 U21826 ( .ip1(\x[32][12] ), .ip2(n17895), .op(n17897) );
  or2_1 U21827 ( .ip1(n24449), .ip2(n17895), .op(n17896) );
  nand2_1 U21828 ( .ip1(n17897), .ip2(n17896), .op(n18497) );
  or2_1 U21829 ( .ip1(n24185), .ip2(\x[32][14] ), .op(n17898) );
  nand2_1 U21830 ( .ip1(n17938), .ip2(n17898), .op(n18505) );
  or2_1 U21831 ( .ip1(n18497), .ip2(n18505), .op(n17935) );
  nor2_1 U21832 ( .ip1(\x[32][13] ), .ip2(n23895), .op(n17899) );
  or2_1 U21833 ( .ip1(n17845), .ip2(n17899), .op(n17902) );
  inv_1 U21834 ( .ip(\x[32][12] ), .op(n17900) );
  or2_1 U21835 ( .ip1(n17900), .ip2(n17899), .op(n17901) );
  nand2_1 U21836 ( .ip1(n17902), .ip2(n17901), .op(n18495) );
  inv_1 U21837 ( .ip(\x[32][11] ), .op(n17929) );
  nor2_1 U21838 ( .ip1(n17929), .ip2(n17981), .op(n17931) );
  buf_1 U21839 ( .ip(n24370), .op(n24451) );
  and2_1 U21840 ( .ip1(n24451), .ip2(\x[32][10] ), .op(n17926) );
  inv_1 U21841 ( .ip(\x[32][9] ), .op(n17924) );
  and2_1 U21842 ( .ip1(n24491), .ip2(\x[32][8] ), .op(n17921) );
  inv_1 U21843 ( .ip(\x[32][6] ), .op(n17919) );
  nor2_1 U21844 ( .ip1(sig_in[6]), .ip2(n17919), .op(n17916) );
  inv_1 U21845 ( .ip(\x[32][4] ), .op(n17914) );
  nor2_1 U21846 ( .ip1(n24462), .ip2(n17914), .op(n17911) );
  inv_1 U21847 ( .ip(\x[32][3] ), .op(n17909) );
  inv_1 U21848 ( .ip(\x[32][1] ), .op(n17904) );
  nor2_1 U21849 ( .ip1(n22513), .ip2(n17904), .op(n17906) );
  inv_1 U21850 ( .ip(\x[32][0] ), .op(n17903) );
  not_ab_or_c_or_d U21851 ( .ip1(n24467), .ip2(n17904), .ip3(sig_in[0]), .ip4(
        n17903), .op(n17905) );
  not_ab_or_c_or_d U21852 ( .ip1(\x[32][2] ), .ip2(n24107), .ip3(n17906), 
        .ip4(n17905), .op(n17908) );
  nor2_1 U21853 ( .ip1(\x[32][2] ), .ip2(n24463), .op(n17907) );
  not_ab_or_c_or_d U21854 ( .ip1(n24251), .ip2(n17909), .ip3(n17908), .ip4(
        n17907), .op(n17910) );
  not_ab_or_c_or_d U21855 ( .ip1(\x[32][3] ), .ip2(n22525), .ip3(n17911), 
        .ip4(n17910), .op(n17913) );
  nor2_1 U21856 ( .ip1(\x[32][5] ), .ip2(n23283), .op(n17912) );
  not_ab_or_c_or_d U21857 ( .ip1(sig_in[4]), .ip2(n17914), .ip3(n17913), .ip4(
        n17912), .op(n17915) );
  not_ab_or_c_or_d U21858 ( .ip1(\x[32][5] ), .ip2(n24482), .ip3(n17916), 
        .ip4(n17915), .op(n17918) );
  nor2_1 U21859 ( .ip1(\x[32][7] ), .ip2(n24492), .op(n17917) );
  not_ab_or_c_or_d U21860 ( .ip1(sig_in[6]), .ip2(n17919), .ip3(n17918), .ip4(
        n17917), .op(n17920) );
  not_ab_or_c_or_d U21861 ( .ip1(\x[32][7] ), .ip2(n24044), .ip3(n17921), 
        .ip4(n17920), .op(n17923) );
  nor2_1 U21862 ( .ip1(\x[32][8] ), .ip2(n23971), .op(n17922) );
  not_ab_or_c_or_d U21863 ( .ip1(sig_in[9]), .ip2(n17924), .ip3(n17923), .ip4(
        n17922), .op(n17925) );
  not_ab_or_c_or_d U21864 ( .ip1(\x[32][9] ), .ip2(n24164), .ip3(n17926), 
        .ip4(n17925), .op(n17928) );
  nor2_1 U21865 ( .ip1(\x[32][10] ), .ip2(n20880), .op(n17927) );
  not_ab_or_c_or_d U21866 ( .ip1(sig_in[11]), .ip2(n17929), .ip3(n17928), 
        .ip4(n17927), .op(n17930) );
  nor2_1 U21867 ( .ip1(n17931), .ip2(n17930), .op(n18496) );
  inv_1 U21868 ( .ip(n18496), .op(n17932) );
  nand2_1 U21869 ( .ip1(n18495), .ip2(n17932), .op(n17933) );
  or2_1 U21870 ( .ip1(n17933), .ip2(n18505), .op(n17934) );
  nand2_1 U21871 ( .ip1(n17935), .ip2(n17934), .op(n17936) );
  not_ab_or_c_or_d U21872 ( .ip1(n17938), .ip2(n18498), .ip3(n17937), .ip4(
        n17936), .op(n24880) );
  nor2_1 U21873 ( .ip1(\x[36][14] ), .ip2(n24327), .op(n17939) );
  or2_1 U21874 ( .ip1(\x[36][15] ), .ip2(n17939), .op(n17941) );
  or2_1 U21875 ( .ip1(n24384), .ip2(n17939), .op(n17940) );
  nand2_1 U21876 ( .ip1(n17941), .ip2(n17940), .op(n18017) );
  or2_1 U21877 ( .ip1(n24081), .ip2(\x[36][13] ), .op(n17942) );
  nand2_1 U21878 ( .ip1(n18017), .ip2(n17942), .op(n18022) );
  or2_1 U21879 ( .ip1(n17845), .ip2(n18022), .op(n17944) );
  inv_1 U21880 ( .ip(\x[36][12] ), .op(n18380) );
  or2_1 U21881 ( .ip1(n18380), .ip2(n18022), .op(n17943) );
  nand2_1 U21882 ( .ip1(n17944), .ip2(n17943), .op(n18420) );
  nand2_1 U21883 ( .ip1(\x[36][11] ), .ip2(n24456), .op(n17974) );
  and2_1 U21884 ( .ip1(n23971), .ip2(\x[36][8] ), .op(n17966) );
  inv_1 U21885 ( .ip(\x[36][7] ), .op(n17964) );
  nor2_1 U21886 ( .ip1(n17732), .ip2(n17964), .op(n17961) );
  inv_1 U21887 ( .ip(\x[36][5] ), .op(n17959) );
  nor2_1 U21888 ( .ip1(n22833), .ip2(n17959), .op(n17956) );
  inv_1 U21889 ( .ip(\x[36][1] ), .op(n17946) );
  inv_1 U21890 ( .ip(\x[36][0] ), .op(n17945) );
  not_ab_or_c_or_d U21891 ( .ip1(n24467), .ip2(n17946), .ip3(sig_in[0]), .ip4(
        n17945), .op(n17950) );
  nand2_1 U21892 ( .ip1(\x[36][1] ), .ip2(n20652), .op(n17948) );
  nand2_1 U21893 ( .ip1(\x[36][3] ), .ip2(n24476), .op(n17947) );
  nand2_1 U21894 ( .ip1(n17948), .ip2(n17947), .op(n17949) );
  not_ab_or_c_or_d U21895 ( .ip1(\x[36][2] ), .ip2(n24335), .ip3(n17950), 
        .ip4(n17949), .op(n17954) );
  nor2_1 U21896 ( .ip1(\x[36][4] ), .ip2(n24256), .op(n17953) );
  nor2_1 U21897 ( .ip1(\x[36][3] ), .ip2(n22795), .op(n17952) );
  not_ab_or_c_or_d U21898 ( .ip1(\x[36][3] ), .ip2(n22795), .ip3(\x[36][2] ), 
        .ip4(n24470), .op(n17951) );
  nor4_1 U21899 ( .ip1(n17954), .ip2(n17953), .ip3(n17952), .ip4(n17951), .op(
        n17955) );
  not_ab_or_c_or_d U21900 ( .ip1(\x[36][4] ), .ip2(n24256), .ip3(n17956), 
        .ip4(n17955), .op(n17958) );
  nor2_1 U21901 ( .ip1(\x[36][6] ), .ip2(n24485), .op(n17957) );
  not_ab_or_c_or_d U21902 ( .ip1(sig_in[5]), .ip2(n17959), .ip3(n17958), .ip4(
        n17957), .op(n17960) );
  not_ab_or_c_or_d U21903 ( .ip1(\x[36][6] ), .ip2(n24355), .ip3(n17961), 
        .ip4(n17960), .op(n17963) );
  nor2_1 U21904 ( .ip1(\x[36][8] ), .ip2(n24358), .op(n17962) );
  not_ab_or_c_or_d U21905 ( .ip1(sig_in[7]), .ip2(n17964), .ip3(n17963), .ip4(
        n17962), .op(n17965) );
  not_ab_or_c_or_d U21906 ( .ip1(\x[36][9] ), .ip2(n23981), .ip3(n17966), 
        .ip4(n17965), .op(n17968) );
  nor2_1 U21907 ( .ip1(\x[36][9] ), .ip2(n24455), .op(n17967) );
  nor2_1 U21908 ( .ip1(n17968), .ip2(n17967), .op(n17969) );
  nand2_1 U21909 ( .ip1(\x[36][10] ), .ip2(n17969), .op(n17972) );
  nor2_1 U21910 ( .ip1(\x[36][11] ), .ip2(n24456), .op(n17971) );
  nor2_1 U21911 ( .ip1(\x[36][10] ), .ip2(n17969), .op(n17970) );
  ab_or_c_or_d U21912 ( .ip1(sig_in[10]), .ip2(n17972), .ip3(n17971), .ip4(
        n17970), .op(n17973) );
  nand2_1 U21913 ( .ip1(n17974), .ip2(n17973), .op(n18381) );
  nor2_1 U21914 ( .ip1(\x[37][13] ), .ip2(n24235), .op(n17975) );
  or2_1 U21915 ( .ip1(n17845), .ip2(n17975), .op(n17978) );
  inv_1 U21916 ( .ip(\x[37][12] ), .op(n17976) );
  or2_1 U21917 ( .ip1(n17976), .ip2(n17975), .op(n17977) );
  nand2_1 U21918 ( .ip1(n17978), .ip2(n17977), .op(n18374) );
  nand2_1 U21919 ( .ip1(n24327), .ip2(\x[37][14] ), .op(n17980) );
  or2_1 U21920 ( .ip1(n24329), .ip2(\x[37][15] ), .op(n18016) );
  nand2_1 U21921 ( .ip1(\x[37][13] ), .ip2(n24235), .op(n17979) );
  nand3_1 U21922 ( .ip1(n17980), .ip2(n18016), .ip3(n17979), .op(n18360) );
  or2_1 U21923 ( .ip1(n18374), .ip2(n18360), .op(n18014) );
  buf_1 U21924 ( .ip(sig_in[11]), .op(n17981) );
  nor2_1 U21925 ( .ip1(n24371), .ip2(\x[37][11] ), .op(n18010) );
  inv_1 U21926 ( .ip(\x[37][9] ), .op(n18006) );
  and2_1 U21927 ( .ip1(n23804), .ip2(\x[37][8] ), .op(n18003) );
  inv_1 U21928 ( .ip(\x[37][4] ), .op(n17993) );
  nor2_1 U21929 ( .ip1(n24462), .ip2(n17993), .op(n17990) );
  inv_1 U21930 ( .ip(\x[37][3] ), .op(n17988) );
  nor2_1 U21931 ( .ip1(\x[37][2] ), .ip2(n24463), .op(n17987) );
  inv_1 U21932 ( .ip(\x[37][1] ), .op(n17983) );
  nor2_1 U21933 ( .ip1(n22513), .ip2(n17983), .op(n17985) );
  inv_1 U21934 ( .ip(\x[37][0] ), .op(n17982) );
  not_ab_or_c_or_d U21935 ( .ip1(n24464), .ip2(n17983), .ip3(sig_in[0]), .ip4(
        n17982), .op(n17984) );
  not_ab_or_c_or_d U21936 ( .ip1(\x[37][2] ), .ip2(n24107), .ip3(n17985), 
        .ip4(n17984), .op(n17986) );
  not_ab_or_c_or_d U21937 ( .ip1(n23251), .ip2(n17988), .ip3(n17987), .ip4(
        n17986), .op(n17989) );
  not_ab_or_c_or_d U21938 ( .ip1(\x[37][3] ), .ip2(n24476), .ip3(n17990), 
        .ip4(n17989), .op(n17992) );
  nor2_1 U21939 ( .ip1(\x[37][5] ), .ip2(n23283), .op(n17991) );
  not_ab_or_c_or_d U21940 ( .ip1(sig_in[4]), .ip2(n17993), .ip3(n17992), .ip4(
        n17991), .op(n17997) );
  nand2_1 U21941 ( .ip1(\x[37][7] ), .ip2(n24492), .op(n17995) );
  nand2_1 U21942 ( .ip1(\x[37][6] ), .ip2(n24485), .op(n17994) );
  nand2_1 U21943 ( .ip1(n17995), .ip2(n17994), .op(n17996) );
  not_ab_or_c_or_d U21944 ( .ip1(\x[37][5] ), .ip2(n24482), .ip3(n17997), 
        .ip4(n17996), .op(n18001) );
  nor2_1 U21945 ( .ip1(\x[37][7] ), .ip2(n24044), .op(n18000) );
  nor2_1 U21946 ( .ip1(\x[37][8] ), .ip2(n24358), .op(n17999) );
  inv_1 U21947 ( .ip(sig_in[6]), .op(n23770) );
  not_ab_or_c_or_d U21948 ( .ip1(\x[37][7] ), .ip2(n24044), .ip3(\x[37][6] ), 
        .ip4(n23770), .op(n17998) );
  nor4_1 U21949 ( .ip1(n18001), .ip2(n18000), .ip3(n17999), .ip4(n17998), .op(
        n18002) );
  not_ab_or_c_or_d U21950 ( .ip1(\x[37][9] ), .ip2(n23981), .ip3(n18003), 
        .ip4(n18002), .op(n18005) );
  nor2_1 U21951 ( .ip1(\x[37][10] ), .ip2(n20880), .op(n18004) );
  not_ab_or_c_or_d U21952 ( .ip1(sig_in[9]), .ip2(n18006), .ip3(n18005), .ip4(
        n18004), .op(n18008) );
  and2_1 U21953 ( .ip1(n24451), .ip2(\x[37][10] ), .op(n18007) );
  not_ab_or_c_or_d U21954 ( .ip1(\x[37][11] ), .ip2(n24136), .ip3(n18008), 
        .ip4(n18007), .op(n18009) );
  nor2_1 U21955 ( .ip1(n18010), .ip2(n18009), .op(n18372) );
  inv_1 U21956 ( .ip(n18372), .op(n18011) );
  nand2_1 U21957 ( .ip1(\x[37][12] ), .ip2(n24233), .op(n18364) );
  nand2_1 U21958 ( .ip1(n18011), .ip2(n18364), .op(n18012) );
  or2_1 U21959 ( .ip1(n18012), .ip2(n18360), .op(n18013) );
  nand2_1 U21960 ( .ip1(n18014), .ip2(n18013), .op(n18026) );
  or2_1 U21961 ( .ip1(n24185), .ip2(\x[37][14] ), .op(n18015) );
  nand2_1 U21962 ( .ip1(\x[37][15] ), .ip2(n24186), .op(n18361) );
  nand2_1 U21963 ( .ip1(n18015), .ip2(n18361), .op(n18371) );
  nand2_1 U21964 ( .ip1(n18371), .ip2(n18016), .op(n18024) );
  nor2_1 U21965 ( .ip1(\x[36][15] ), .ip2(n24090), .op(n18384) );
  or2_1 U21966 ( .ip1(n18017), .ip2(n18384), .op(n18021) );
  nand2_1 U21967 ( .ip1(\x[36][13] ), .ip2(n24235), .op(n18019) );
  nand2_1 U21968 ( .ip1(\x[36][14] ), .ip2(n23938), .op(n18018) );
  nand2_1 U21969 ( .ip1(n18019), .ip2(n18018), .op(n18382) );
  or2_1 U21970 ( .ip1(n18382), .ip2(n18384), .op(n18020) );
  nand2_1 U21971 ( .ip1(n18021), .ip2(n18020), .op(n18422) );
  or3_1 U21972 ( .ip1(n18022), .ip2(n18380), .ip3(n17845), .op(n18023) );
  nand3_1 U21973 ( .ip1(n18024), .ip2(n18422), .ip3(n18023), .op(n18025) );
  not_ab_or_c_or_d U21974 ( .ip1(n18420), .ip2(n18381), .ip3(n18026), .ip4(
        n18025), .op(n24874) );
  and2_1 U21975 ( .ip1(n23895), .ip2(\x[38][13] ), .op(n18027) );
  nor2_1 U21976 ( .ip1(\x[38][15] ), .ip2(n24090), .op(n18032) );
  not_ab_or_c_or_d U21977 ( .ip1(\x[38][14] ), .ip2(n24185), .ip3(n18027), 
        .ip4(n18032), .op(n18370) );
  nand2_1 U21978 ( .ip1(\x[38][12] ), .ip2(n24233), .op(n18028) );
  nand2_1 U21979 ( .ip1(n18370), .ip2(n18028), .op(n18358) );
  nor2_1 U21980 ( .ip1(\x[38][14] ), .ip2(n24327), .op(n18029) );
  or2_1 U21981 ( .ip1(\x[38][15] ), .ip2(n18029), .op(n18031) );
  or2_1 U21982 ( .ip1(n24329), .ip2(n18029), .op(n18030) );
  nand2_1 U21983 ( .ip1(n18031), .ip2(n18030), .op(n18074) );
  nor2_1 U21984 ( .ip1(n18032), .ip2(n18074), .op(n18368) );
  inv_1 U21985 ( .ip(n18368), .op(n18124) );
  nor2_1 U21986 ( .ip1(\x[38][13] ), .ip2(n24332), .op(n18033) );
  or2_1 U21987 ( .ip1(sig_in[12]), .ip2(n18033), .op(n18036) );
  inv_1 U21988 ( .ip(\x[38][12] ), .op(n18034) );
  or2_1 U21989 ( .ip1(n18034), .ip2(n18033), .op(n18035) );
  nand2_1 U21990 ( .ip1(n18036), .ip2(n18035), .op(n18359) );
  nor2_1 U21991 ( .ip1(\x[38][11] ), .ip2(n24456), .op(n18073) );
  and2_1 U21992 ( .ip1(n24451), .ip2(\x[38][10] ), .op(n18071) );
  inv_1 U21993 ( .ip(\x[38][9] ), .op(n18068) );
  and2_1 U21994 ( .ip1(n24100), .ip2(\x[38][8] ), .op(n18065) );
  inv_1 U21995 ( .ip(\x[38][7] ), .op(n18063) );
  inv_1 U21996 ( .ip(\x[38][6] ), .op(n18055) );
  nor2_1 U21997 ( .ip1(sig_in[6]), .ip2(n18055), .op(n18053) );
  nor2_1 U21998 ( .ip1(n24347), .ip2(\x[38][4] ), .op(n18047) );
  inv_1 U21999 ( .ip(\x[38][3] ), .op(n18043) );
  nor2_1 U22000 ( .ip1(sig_in[3]), .ip2(n18043), .op(n18045) );
  inv_1 U22001 ( .ip(\x[38][1] ), .op(n18038) );
  nor2_1 U22002 ( .ip1(n22513), .ip2(n18038), .op(n18040) );
  inv_1 U22003 ( .ip(\x[38][0] ), .op(n18037) );
  not_ab_or_c_or_d U22004 ( .ip1(n24467), .ip2(n18038), .ip3(sig_in[0]), .ip4(
        n18037), .op(n18039) );
  not_ab_or_c_or_d U22005 ( .ip1(\x[38][2] ), .ip2(n24335), .ip3(n18040), 
        .ip4(n18039), .op(n18042) );
  nor2_1 U22006 ( .ip1(\x[38][2] ), .ip2(n24463), .op(n18041) );
  not_ab_or_c_or_d U22007 ( .ip1(n23251), .ip2(n18043), .ip3(n18042), .ip4(
        n18041), .op(n18044) );
  not_ab_or_c_or_d U22008 ( .ip1(\x[38][4] ), .ip2(n23860), .ip3(n18045), 
        .ip4(n18044), .op(n18046) );
  or2_1 U22009 ( .ip1(n18047), .ip2(n18046), .op(n18048) );
  or2_1 U22010 ( .ip1(sig_in[5]), .ip2(n18048), .op(n18051) );
  inv_1 U22011 ( .ip(\x[38][5] ), .op(n18049) );
  or2_1 U22012 ( .ip1(n18049), .ip2(n18048), .op(n18050) );
  nand2_1 U22013 ( .ip1(n18051), .ip2(n18050), .op(n18052) );
  not_ab_or_c_or_d U22014 ( .ip1(\x[38][5] ), .ip2(n24482), .ip3(n18053), 
        .ip4(n18052), .op(n18054) );
  or2_1 U22015 ( .ip1(sig_in[6]), .ip2(n18054), .op(n18057) );
  or2_1 U22016 ( .ip1(n18055), .ip2(n18054), .op(n18056) );
  nand2_1 U22017 ( .ip1(n18057), .ip2(n18056), .op(n18058) );
  or2_1 U22018 ( .ip1(\x[38][7] ), .ip2(n18058), .op(n18060) );
  or2_1 U22019 ( .ip1(n24044), .ip2(n18058), .op(n18059) );
  nand2_1 U22020 ( .ip1(n18060), .ip2(n18059), .op(n18062) );
  nor2_1 U22021 ( .ip1(\x[38][8] ), .ip2(n23971), .op(n18061) );
  not_ab_or_c_or_d U22022 ( .ip1(sig_in[7]), .ip2(n18063), .ip3(n18062), .ip4(
        n18061), .op(n18064) );
  not_ab_or_c_or_d U22023 ( .ip1(\x[38][9] ), .ip2(n24164), .ip3(n18065), 
        .ip4(n18064), .op(n18067) );
  nor2_1 U22024 ( .ip1(\x[38][10] ), .ip2(n20880), .op(n18066) );
  not_ab_or_c_or_d U22025 ( .ip1(sig_in[9]), .ip2(n18068), .ip3(n18067), .ip4(
        n18066), .op(n18070) );
  inv_1 U22026 ( .ip(n17981), .op(n24239) );
  and2_1 U22027 ( .ip1(n24239), .ip2(\x[38][11] ), .op(n18069) );
  nor3_1 U22028 ( .ip1(n18071), .ip2(n18070), .ip3(n18069), .op(n18072) );
  nor2_1 U22029 ( .ip1(n18073), .ip2(n18072), .op(n18357) );
  and3_1 U22030 ( .ip1(n18074), .ip2(n18359), .ip3(n18357), .op(n18123) );
  and2_1 U22031 ( .ip1(n24332), .ip2(\x[39][13] ), .op(n18075) );
  or2_1 U22032 ( .ip1(\x[39][12] ), .ip2(n18075), .op(n18077) );
  or2_1 U22033 ( .ip1(n24079), .ip2(n18075), .op(n18076) );
  nand2_1 U22034 ( .ip1(n18077), .ip2(n18076), .op(n18338) );
  nor2_1 U22035 ( .ip1(\x[39][10] ), .ip2(n20880), .op(n18111) );
  nor2_1 U22036 ( .ip1(n17981), .ip2(n18111), .op(n18078) );
  nor2_1 U22037 ( .ip1(\x[39][11] ), .ip2(n18078), .op(n18110) );
  inv_1 U22038 ( .ip(\x[39][7] ), .op(n18100) );
  and2_1 U22039 ( .ip1(n24335), .ip2(\x[39][2] ), .op(n18087) );
  inv_1 U22040 ( .ip(\x[39][1] ), .op(n18080) );
  inv_1 U22041 ( .ip(\x[39][0] ), .op(n18079) );
  not_ab_or_c_or_d U22042 ( .ip1(n24464), .ip2(n18080), .ip3(sig_in[0]), .ip4(
        n18079), .op(n18081) );
  or2_1 U22043 ( .ip1(\x[39][1] ), .ip2(n18081), .op(n18083) );
  or2_1 U22044 ( .ip1(n21685), .ip2(n18081), .op(n18082) );
  nand2_1 U22045 ( .ip1(n18083), .ip2(n18082), .op(n18085) );
  nor2_1 U22046 ( .ip1(\x[39][2] ), .ip2(n24463), .op(n18084) );
  nor2_1 U22047 ( .ip1(n18085), .ip2(n18084), .op(n18086) );
  not_ab_or_c_or_d U22048 ( .ip1(\x[39][3] ), .ip2(n22795), .ip3(n18087), 
        .ip4(n18086), .op(n18090) );
  nor2_1 U22049 ( .ip1(\x[39][5] ), .ip2(n23283), .op(n18091) );
  nor2_1 U22050 ( .ip1(\x[39][3] ), .ip2(n24342), .op(n18089) );
  nor2_1 U22051 ( .ip1(\x[39][4] ), .ip2(n24256), .op(n18088) );
  nor4_1 U22052 ( .ip1(n18090), .ip2(n18091), .ip3(n18089), .ip4(n18088), .op(
        n18097) );
  nand2_1 U22053 ( .ip1(n23770), .ip2(\x[39][6] ), .op(n18095) );
  inv_1 U22054 ( .ip(n18091), .op(n18092) );
  nand3_1 U22055 ( .ip1(\x[39][4] ), .ip2(n23721), .ip3(n18092), .op(n18094)
         );
  nand2_1 U22056 ( .ip1(\x[39][7] ), .ip2(n24461), .op(n18093) );
  nand3_1 U22057 ( .ip1(n18095), .ip2(n18094), .ip3(n18093), .op(n18096) );
  not_ab_or_c_or_d U22058 ( .ip1(\x[39][5] ), .ip2(n24482), .ip3(n18097), 
        .ip4(n18096), .op(n18099) );
  not_ab_or_c_or_d U22059 ( .ip1(\x[39][7] ), .ip2(n24142), .ip3(\x[39][6] ), 
        .ip4(n23770), .op(n18098) );
  not_ab_or_c_or_d U22060 ( .ip1(sig_in[7]), .ip2(n18100), .ip3(n18099), .ip4(
        n18098), .op(n18101) );
  nand2_1 U22061 ( .ip1(\x[39][8] ), .ip2(n18101), .op(n18104) );
  inv_1 U22062 ( .ip(n21171), .op(n24269) );
  nor2_1 U22063 ( .ip1(\x[39][9] ), .ip2(n24269), .op(n18103) );
  nor2_1 U22064 ( .ip1(\x[39][8] ), .ip2(n18101), .op(n18102) );
  ab_or_c_or_d U22065 ( .ip1(n23779), .ip2(n18104), .ip3(n18103), .ip4(n18102), 
        .op(n18108) );
  nand2_1 U22066 ( .ip1(\x[39][9] ), .ip2(n24164), .op(n18107) );
  nand2_1 U22067 ( .ip1(\x[39][11] ), .ip2(n24456), .op(n18106) );
  nand2_1 U22068 ( .ip1(\x[39][10] ), .ip2(n23980), .op(n18105) );
  and4_1 U22069 ( .ip1(n18108), .ip2(n18107), .ip3(n18106), .ip4(n18105), .op(
        n18109) );
  ab_or_c_or_d U22070 ( .ip1(n18111), .ip2(n17981), .ip3(n18110), .ip4(n18109), 
        .op(n18334) );
  nand2_1 U22071 ( .ip1(n18338), .ip2(n18334), .op(n18113) );
  nor2_1 U22072 ( .ip1(\x[39][12] ), .ip2(n24233), .op(n18333) );
  nor2_1 U22073 ( .ip1(\x[39][13] ), .ip2(n24137), .op(n18336) );
  nor2_1 U22074 ( .ip1(n18333), .ip2(n18336), .op(n18112) );
  nand2_1 U22075 ( .ip1(n18113), .ip2(n18112), .op(n18116) );
  nor2_1 U22076 ( .ip1(\x[39][15] ), .ip2(n24090), .op(n18117) );
  or2_1 U22077 ( .ip1(\x[39][14] ), .ip2(n18117), .op(n18115) );
  or2_1 U22078 ( .ip1(n24185), .ip2(n18117), .op(n18114) );
  nand2_1 U22079 ( .ip1(n18115), .ip2(n18114), .op(n18341) );
  nand2_1 U22080 ( .ip1(n18116), .ip2(n18341), .op(n18121) );
  inv_1 U22081 ( .ip(n18117), .op(n18119) );
  nand2_1 U22082 ( .ip1(\x[39][15] ), .ip2(n24186), .op(n18339) );
  or2_1 U22083 ( .ip1(n24185), .ip2(\x[39][14] ), .op(n18118) );
  nand2_1 U22084 ( .ip1(n18339), .ip2(n18118), .op(n18335) );
  nand2_1 U22085 ( .ip1(n18119), .ip2(n18335), .op(n18120) );
  nand2_1 U22086 ( .ip1(n18121), .ip2(n18120), .op(n18122) );
  not_ab_or_c_or_d U22087 ( .ip1(n18358), .ip2(n18124), .ip3(n18123), .ip4(
        n18122), .op(n24862) );
  nor2_1 U22088 ( .ip1(\x[40][15] ), .ip2(n24090), .op(n18342) );
  nor2_1 U22089 ( .ip1(\x[40][13] ), .ip2(n24235), .op(n18125) );
  or2_1 U22090 ( .ip1(n17845), .ip2(n18125), .op(n18128) );
  inv_1 U22091 ( .ip(\x[40][12] ), .op(n18126) );
  or2_1 U22092 ( .ip1(n18126), .ip2(n18125), .op(n18127) );
  nand2_1 U22093 ( .ip1(n18128), .ip2(n18127), .op(n18346) );
  and2_1 U22094 ( .ip1(n24451), .ip2(\x[40][10] ), .op(n18155) );
  and2_1 U22095 ( .ip1(n24043), .ip2(\x[40][9] ), .op(n18149) );
  and2_1 U22096 ( .ip1(n24461), .ip2(\x[40][7] ), .op(n18145) );
  inv_1 U22097 ( .ip(\x[40][3] ), .op(n18135) );
  nor2_1 U22098 ( .ip1(\x[40][2] ), .ip2(n24463), .op(n18134) );
  inv_1 U22099 ( .ip(\x[40][1] ), .op(n18130) );
  nor2_1 U22100 ( .ip1(n22513), .ip2(n18130), .op(n18132) );
  inv_1 U22101 ( .ip(\x[40][0] ), .op(n18129) );
  not_ab_or_c_or_d U22102 ( .ip1(sig_in[1]), .ip2(n18130), .ip3(sig_in[0]), 
        .ip4(n18129), .op(n18131) );
  not_ab_or_c_or_d U22103 ( .ip1(\x[40][2] ), .ip2(n24107), .ip3(n18132), 
        .ip4(n18131), .op(n18133) );
  not_ab_or_c_or_d U22104 ( .ip1(n24251), .ip2(n18135), .ip3(n18134), .ip4(
        n18133), .op(n18139) );
  nand2_1 U22105 ( .ip1(\x[40][5] ), .ip2(n24119), .op(n18137) );
  nand2_1 U22106 ( .ip1(\x[40][4] ), .ip2(n24347), .op(n18136) );
  nand2_1 U22107 ( .ip1(n18137), .ip2(n18136), .op(n18138) );
  not_ab_or_c_or_d U22108 ( .ip1(\x[40][3] ), .ip2(n22795), .ip3(n18139), 
        .ip4(n18138), .op(n18143) );
  inv_1 U22109 ( .ip(sig_in[6]), .op(n24355) );
  nor2_1 U22110 ( .ip1(\x[40][6] ), .ip2(n24355), .op(n18142) );
  nor2_1 U22111 ( .ip1(\x[40][5] ), .ip2(n23283), .op(n18141) );
  not_ab_or_c_or_d U22112 ( .ip1(\x[40][5] ), .ip2(n24482), .ip3(\x[40][4] ), 
        .ip4(n24347), .op(n18140) );
  nor4_1 U22113 ( .ip1(n18143), .ip2(n18142), .ip3(n18141), .ip4(n18140), .op(
        n18144) );
  not_ab_or_c_or_d U22114 ( .ip1(\x[40][6] ), .ip2(n23770), .ip3(n18145), 
        .ip4(n18144), .op(n18147) );
  nor2_1 U22115 ( .ip1(\x[40][7] ), .ip2(n24142), .op(n18146) );
  nor2_1 U22116 ( .ip1(n18147), .ip2(n18146), .op(n18148) );
  not_ab_or_c_or_d U22117 ( .ip1(\x[40][8] ), .ip2(n24491), .ip3(n18149), 
        .ip4(n18148), .op(n18153) );
  not_ab_or_c_or_d U22118 ( .ip1(\x[40][9] ), .ip2(n24043), .ip3(\x[40][8] ), 
        .ip4(n24358), .op(n18152) );
  nor2_1 U22119 ( .ip1(\x[40][10] ), .ip2(n20880), .op(n18151) );
  nor2_1 U22120 ( .ip1(\x[40][9] ), .ip2(n24269), .op(n18150) );
  nor4_1 U22121 ( .ip1(n18153), .ip2(n18152), .ip3(n18151), .ip4(n18150), .op(
        n18154) );
  not_ab_or_c_or_d U22122 ( .ip1(\x[40][11] ), .ip2(n24136), .ip3(n18155), 
        .ip4(n18154), .op(n18157) );
  nor2_1 U22123 ( .ip1(\x[40][11] ), .ip2(n24456), .op(n18156) );
  nor2_1 U22124 ( .ip1(n18157), .ip2(n18156), .op(n18347) );
  nand2_1 U22125 ( .ip1(n24230), .ip2(\x[40][14] ), .op(n18344) );
  inv_1 U22126 ( .ip(n18344), .op(n18160) );
  nand2_1 U22127 ( .ip1(\x[40][13] ), .ip2(n24235), .op(n18159) );
  inv_1 U22128 ( .ip(n17845), .op(n24450) );
  nand2_1 U22129 ( .ip1(\x[40][12] ), .ip2(n24450), .op(n18158) );
  nand2_1 U22130 ( .ip1(n18159), .ip2(n18158), .op(n18348) );
  not_ab_or_c_or_d U22131 ( .ip1(n18346), .ip2(n18347), .ip3(n18160), .ip4(
        n18348), .op(n18163) );
  or2_1 U22132 ( .ip1(n24185), .ip2(\x[40][14] ), .op(n18162) );
  nand2_1 U22133 ( .ip1(\x[40][15] ), .ip2(n24186), .op(n18161) );
  nand2_1 U22134 ( .ip1(n18162), .ip2(n18161), .op(n18343) );
  nor2_1 U22135 ( .ip1(n18163), .ip2(n18343), .op(n18212) );
  nor2_1 U22136 ( .ip1(\x[41][15] ), .ip2(n24090), .op(n18168) );
  buf_1 U22137 ( .ip(n24329), .op(n23143) );
  nand2_1 U22138 ( .ip1(n23143), .ip2(\x[41][15] ), .op(n18308) );
  inv_1 U22139 ( .ip(n18308), .op(n18164) );
  or2_1 U22140 ( .ip1(sig_in[14]), .ip2(n18164), .op(n18167) );
  inv_1 U22141 ( .ip(\x[41][14] ), .op(n18165) );
  or2_1 U22142 ( .ip1(n18165), .ip2(n18164), .op(n18166) );
  nand2_1 U22143 ( .ip1(n18167), .ip2(n18166), .op(n18328) );
  nor2_1 U22144 ( .ip1(n18168), .ip2(n18328), .op(n18211) );
  and2_1 U22145 ( .ip1(n24235), .ip2(\x[41][13] ), .op(n18169) );
  not_ab_or_c_or_d U22146 ( .ip1(\x[41][14] ), .ip2(n24185), .ip3(n18169), 
        .ip4(n18168), .op(n18306) );
  nor2_1 U22147 ( .ip1(\x[41][13] ), .ip2(n24376), .op(n18171) );
  nor2_1 U22148 ( .ip1(\x[41][12] ), .ip2(n24233), .op(n18170) );
  nor2_1 U22149 ( .ip1(n18171), .ip2(n18170), .op(n18329) );
  inv_1 U22150 ( .ip(n18329), .op(n18172) );
  nand2_1 U22151 ( .ip1(n18306), .ip2(n18172), .op(n18209) );
  nand2_1 U22152 ( .ip1(\x[41][12] ), .ip2(n24233), .op(n18305) );
  inv_1 U22153 ( .ip(\x[41][11] ), .op(n18204) );
  and2_1 U22154 ( .ip1(n24451), .ip2(\x[41][10] ), .op(n18201) );
  nor2_1 U22155 ( .ip1(\x[41][7] ), .ip2(n24142), .op(n18192) );
  inv_1 U22156 ( .ip(\x[41][6] ), .op(n18173) );
  nor3_1 U22157 ( .ip1(sig_in[6]), .ip2(n18192), .ip3(n18173), .op(n18195) );
  and2_1 U22158 ( .ip1(n23283), .ip2(\x[41][5] ), .op(n18189) );
  inv_1 U22159 ( .ip(\x[41][3] ), .op(n18180) );
  inv_1 U22160 ( .ip(\x[41][1] ), .op(n18175) );
  nor2_1 U22161 ( .ip1(n24467), .ip2(n18175), .op(n18177) );
  inv_1 U22162 ( .ip(\x[41][0] ), .op(n18174) );
  not_ab_or_c_or_d U22163 ( .ip1(n24467), .ip2(n18175), .ip3(sig_in[0]), .ip4(
        n18174), .op(n18176) );
  not_ab_or_c_or_d U22164 ( .ip1(\x[41][2] ), .ip2(n24335), .ip3(n18177), 
        .ip4(n18176), .op(n18179) );
  nor2_1 U22165 ( .ip1(\x[41][2] ), .ip2(n24463), .op(n18178) );
  not_ab_or_c_or_d U22166 ( .ip1(n23251), .ip2(n18180), .ip3(n18179), .ip4(
        n18178), .op(n18181) );
  or2_1 U22167 ( .ip1(\x[41][3] ), .ip2(n18181), .op(n18183) );
  or2_1 U22168 ( .ip1(n22525), .ip2(n18181), .op(n18182) );
  nand2_1 U22169 ( .ip1(n18183), .ip2(n18182), .op(n18184) );
  or2_1 U22170 ( .ip1(sig_in[4]), .ip2(n18184), .op(n18187) );
  inv_1 U22171 ( .ip(\x[41][4] ), .op(n18185) );
  or2_1 U22172 ( .ip1(n18185), .ip2(n18184), .op(n18186) );
  nand2_1 U22173 ( .ip1(n18187), .ip2(n18186), .op(n18188) );
  not_ab_or_c_or_d U22174 ( .ip1(\x[41][4] ), .ip2(n23860), .ip3(n18189), 
        .ip4(n18188), .op(n18193) );
  nor2_1 U22175 ( .ip1(\x[41][6] ), .ip2(n24485), .op(n18191) );
  nor2_1 U22176 ( .ip1(\x[41][5] ), .ip2(n23283), .op(n18190) );
  nor4_1 U22177 ( .ip1(n18193), .ip2(n18192), .ip3(n18191), .ip4(n18190), .op(
        n18194) );
  not_ab_or_c_or_d U22178 ( .ip1(\x[41][7] ), .ip2(n24492), .ip3(n18195), 
        .ip4(n18194), .op(n18199) );
  nand2_1 U22179 ( .ip1(\x[41][8] ), .ip2(n24100), .op(n18198) );
  nor2_1 U22180 ( .ip1(\x[41][8] ), .ip2(n23971), .op(n18197) );
  nor2_1 U22181 ( .ip1(\x[41][9] ), .ip2(n24455), .op(n18196) );
  not_ab_or_c_or_d U22182 ( .ip1(n18199), .ip2(n18198), .ip3(n18197), .ip4(
        n18196), .op(n18200) );
  not_ab_or_c_or_d U22183 ( .ip1(\x[41][9] ), .ip2(n24269), .ip3(n18201), 
        .ip4(n18200), .op(n18203) );
  nor2_1 U22184 ( .ip1(\x[41][10] ), .ip2(n20880), .op(n18202) );
  not_ab_or_c_or_d U22185 ( .ip1(sig_in[11]), .ip2(n18204), .ip3(n18203), 
        .ip4(n18202), .op(n18205) );
  or2_1 U22186 ( .ip1(\x[41][11] ), .ip2(n18205), .op(n18207) );
  or2_1 U22187 ( .ip1(n24136), .ip2(n18205), .op(n18206) );
  nand2_1 U22188 ( .ip1(n18207), .ip2(n18206), .op(n18326) );
  nand3_1 U22189 ( .ip1(n18306), .ip2(n18305), .ip3(n18326), .op(n18208) );
  nand2_1 U22190 ( .ip1(n18209), .ip2(n18208), .op(n18210) );
  nor4_1 U22191 ( .ip1(n18342), .ip2(n18212), .ip3(n18211), .ip4(n18210), .op(
        n24859) );
  nand2_1 U22192 ( .ip1(\x[42][15] ), .ip2(n24186), .op(n18255) );
  and2_1 U22193 ( .ip1(\x[42][14] ), .ip2(n24230), .op(n18213) );
  nor2_1 U22194 ( .ip1(n24384), .ip2(\x[42][15] ), .op(n18309) );
  nor2_1 U22195 ( .ip1(n18213), .ip2(n18309), .op(n18325) );
  inv_1 U22196 ( .ip(n18325), .op(n18319) );
  nor2_1 U22197 ( .ip1(\x[43][15] ), .ip2(n23143), .op(n18294) );
  nor2_1 U22198 ( .ip1(\x[43][14] ), .ip2(n24327), .op(n18214) );
  or2_1 U22199 ( .ip1(\x[43][15] ), .ip2(n18214), .op(n18216) );
  or2_1 U22200 ( .ip1(n24180), .ip2(n18214), .op(n18215) );
  nand2_1 U22201 ( .ip1(n18216), .ip2(n18215), .op(n19378) );
  nor2_1 U22202 ( .ip1(n18294), .ip2(n19378), .op(n18254) );
  and2_1 U22203 ( .ip1(\x[42][11] ), .ip2(n24239), .op(n18219) );
  nor2_1 U22204 ( .ip1(\x[42][11] ), .ip2(n24456), .op(n18218) );
  nor2_1 U22205 ( .ip1(\x[42][10] ), .ip2(n20880), .op(n18217) );
  nor2_1 U22206 ( .ip1(n18218), .ip2(n18217), .op(n18247) );
  or2_1 U22207 ( .ip1(n18219), .ip2(n18247), .op(n18321) );
  and2_1 U22208 ( .ip1(n24451), .ip2(\x[42][10] ), .op(n18220) );
  not_ab_or_c_or_d U22209 ( .ip1(\x[42][9] ), .ip2(n24043), .ip3(n18220), 
        .ip4(n18219), .op(n18316) );
  inv_1 U22210 ( .ip(\x[42][8] ), .op(n18244) );
  nor2_1 U22211 ( .ip1(n24455), .ip2(\x[42][9] ), .op(n18243) );
  or3_1 U22212 ( .ip1(n23779), .ip2(n18244), .ip3(n18243), .op(n18221) );
  nand2_1 U22213 ( .ip1(n18316), .ip2(n18221), .op(n18222) );
  nand2_1 U22214 ( .ip1(n18321), .ip2(n18222), .op(n18252) );
  inv_1 U22215 ( .ip(\x[42][7] ), .op(n18240) );
  nor2_1 U22216 ( .ip1(n17732), .ip2(n18240), .op(n18238) );
  inv_1 U22217 ( .ip(\x[42][5] ), .op(n18236) );
  nor2_1 U22218 ( .ip1(n22833), .ip2(n18236), .op(n18233) );
  inv_1 U22219 ( .ip(\x[42][3] ), .op(n18231) );
  inv_1 U22220 ( .ip(sig_in[3]), .op(n22795) );
  and2_1 U22221 ( .ip1(n24335), .ip2(\x[42][2] ), .op(n18228) );
  nand2_1 U22222 ( .ip1(\x[42][1] ), .ip2(n21685), .op(n18226) );
  nand2_1 U22223 ( .ip1(\x[42][0] ), .ip2(n24143), .op(n18225) );
  nor2_1 U22224 ( .ip1(\x[42][2] ), .ip2(n24463), .op(n18224) );
  nor2_1 U22225 ( .ip1(\x[42][1] ), .ip2(n21685), .op(n18223) );
  not_ab_or_c_or_d U22226 ( .ip1(n18226), .ip2(n18225), .ip3(n18224), .ip4(
        n18223), .op(n18227) );
  not_ab_or_c_or_d U22227 ( .ip1(\x[42][3] ), .ip2(n22795), .ip3(n18228), 
        .ip4(n18227), .op(n18230) );
  nor2_1 U22228 ( .ip1(\x[42][4] ), .ip2(n24256), .op(n18229) );
  not_ab_or_c_or_d U22229 ( .ip1(n24251), .ip2(n18231), .ip3(n18230), .ip4(
        n18229), .op(n18232) );
  not_ab_or_c_or_d U22230 ( .ip1(\x[42][4] ), .ip2(n24347), .ip3(n18233), 
        .ip4(n18232), .op(n18235) );
  nor2_1 U22231 ( .ip1(\x[42][6] ), .ip2(n24355), .op(n18234) );
  not_ab_or_c_or_d U22232 ( .ip1(n22833), .ip2(n18236), .ip3(n18235), .ip4(
        n18234), .op(n18237) );
  not_ab_or_c_or_d U22233 ( .ip1(\x[42][6] ), .ip2(n23509), .ip3(n18238), 
        .ip4(n18237), .op(n18239) );
  or2_1 U22234 ( .ip1(sig_in[7]), .ip2(n18239), .op(n18242) );
  or2_1 U22235 ( .ip1(n18240), .ip2(n18239), .op(n18241) );
  nand2_1 U22236 ( .ip1(n18242), .ip2(n18241), .op(n18311) );
  or2_1 U22237 ( .ip1(sig_in[8]), .ip2(n18243), .op(n18246) );
  or2_1 U22238 ( .ip1(n18244), .ip2(n18243), .op(n18245) );
  nand2_1 U22239 ( .ip1(n18246), .ip2(n18245), .op(n18314) );
  nand3_1 U22240 ( .ip1(n18247), .ip2(n18311), .ip3(n18314), .op(n18251) );
  or2_1 U22241 ( .ip1(n24185), .ip2(\x[42][14] ), .op(n18248) );
  nand2_1 U22242 ( .ip1(n18255), .ip2(n18248), .op(n18298) );
  nor2_1 U22243 ( .ip1(\x[42][13] ), .ip2(n24081), .op(n18250) );
  nor2_1 U22244 ( .ip1(\x[42][12] ), .ip2(n24233), .op(n18249) );
  or2_1 U22245 ( .ip1(n18250), .ip2(n18249), .op(n18324) );
  not_ab_or_c_or_d U22246 ( .ip1(n18252), .ip2(n18251), .ip3(n18298), .ip4(
        n18324), .op(n18253) );
  not_ab_or_c_or_d U22247 ( .ip1(n18255), .ip2(n18319), .ip3(n18254), .ip4(
        n18253), .op(n18304) );
  inv_1 U22248 ( .ip(n21171), .op(n24164) );
  nor2_1 U22249 ( .ip1(\x[43][9] ), .ip2(n24164), .op(n18280) );
  inv_1 U22250 ( .ip(\x[43][8] ), .op(n18256) );
  nor3_1 U22251 ( .ip1(sig_in[8]), .ip2(n18280), .ip3(n18256), .op(n18283) );
  and2_1 U22252 ( .ip1(n24461), .ip2(\x[43][7] ), .op(n18277) );
  inv_1 U22253 ( .ip(\x[43][5] ), .op(n18275) );
  inv_1 U22254 ( .ip(\x[43][4] ), .op(n18267) );
  nor2_1 U22255 ( .ip1(n24462), .ip2(n18267), .op(n18265) );
  inv_1 U22256 ( .ip(\x[43][3] ), .op(n18263) );
  inv_1 U22257 ( .ip(\x[43][1] ), .op(n18258) );
  nor2_1 U22258 ( .ip1(n22513), .ip2(n18258), .op(n18260) );
  inv_1 U22259 ( .ip(\x[43][0] ), .op(n18257) );
  not_ab_or_c_or_d U22260 ( .ip1(n24467), .ip2(n18258), .ip3(sig_in[0]), .ip4(
        n18257), .op(n18259) );
  not_ab_or_c_or_d U22261 ( .ip1(\x[43][2] ), .ip2(n24107), .ip3(n18260), 
        .ip4(n18259), .op(n18262) );
  nor2_1 U22262 ( .ip1(\x[43][2] ), .ip2(n24463), .op(n18261) );
  not_ab_or_c_or_d U22263 ( .ip1(n24251), .ip2(n18263), .ip3(n18262), .ip4(
        n18261), .op(n18264) );
  not_ab_or_c_or_d U22264 ( .ip1(\x[43][3] ), .ip2(n22795), .ip3(n18265), 
        .ip4(n18264), .op(n18266) );
  or2_1 U22265 ( .ip1(sig_in[4]), .ip2(n18266), .op(n18269) );
  or2_1 U22266 ( .ip1(n18267), .ip2(n18266), .op(n18268) );
  nand2_1 U22267 ( .ip1(n18269), .ip2(n18268), .op(n18270) );
  or2_1 U22268 ( .ip1(\x[43][5] ), .ip2(n18270), .op(n18272) );
  or2_1 U22269 ( .ip1(n24482), .ip2(n18270), .op(n18271) );
  nand2_1 U22270 ( .ip1(n18272), .ip2(n18271), .op(n18274) );
  nor2_1 U22271 ( .ip1(\x[43][6] ), .ip2(n23509), .op(n18273) );
  not_ab_or_c_or_d U22272 ( .ip1(sig_in[5]), .ip2(n18275), .ip3(n18274), .ip4(
        n18273), .op(n18276) );
  not_ab_or_c_or_d U22273 ( .ip1(\x[43][6] ), .ip2(n24355), .ip3(n18277), 
        .ip4(n18276), .op(n18281) );
  nor2_1 U22274 ( .ip1(\x[43][7] ), .ip2(n24142), .op(n18279) );
  nor2_1 U22275 ( .ip1(\x[43][8] ), .ip2(n23971), .op(n18278) );
  nor4_1 U22276 ( .ip1(n18281), .ip2(n18280), .ip3(n18279), .ip4(n18278), .op(
        n18282) );
  not_ab_or_c_or_d U22277 ( .ip1(\x[43][9] ), .ip2(n24164), .ip3(n18283), 
        .ip4(n18282), .op(n18287) );
  nand2_1 U22278 ( .ip1(\x[43][10] ), .ip2(n24370), .op(n18286) );
  nor2_1 U22279 ( .ip1(\x[43][10] ), .ip2(n20880), .op(n18285) );
  nor2_1 U22280 ( .ip1(\x[43][11] ), .ip2(n21793), .op(n18284) );
  not_ab_or_c_or_d U22281 ( .ip1(n18287), .ip2(n18286), .ip3(n18285), .ip4(
        n18284), .op(n18288) );
  or2_1 U22282 ( .ip1(\x[43][11] ), .ip2(n18288), .op(n18290) );
  or2_1 U22283 ( .ip1(n24136), .ip2(n18288), .op(n18289) );
  nand2_1 U22284 ( .ip1(n18290), .ip2(n18289), .op(n19319) );
  and2_1 U22285 ( .ip1(n24235), .ip2(\x[43][13] ), .op(n18291) );
  or2_1 U22286 ( .ip1(\x[43][12] ), .ip2(n18291), .op(n18293) );
  or2_1 U22287 ( .ip1(n24079), .ip2(n18291), .op(n18292) );
  nand2_1 U22288 ( .ip1(n18293), .ip2(n18292), .op(n19322) );
  inv_1 U22289 ( .ip(n18294), .op(n19373) );
  nand2_1 U22290 ( .ip1(n23938), .ip2(\x[43][14] ), .op(n19321) );
  and2_1 U22291 ( .ip1(n19373), .ip2(n19321), .op(n18297) );
  nand3_1 U22292 ( .ip1(n19319), .ip2(n19322), .ip3(n18297), .op(n18303) );
  nor2_1 U22293 ( .ip1(\x[43][13] ), .ip2(n23895), .op(n18296) );
  nor2_1 U22294 ( .ip1(\x[43][12] ), .ip2(n24450), .op(n18295) );
  or2_1 U22295 ( .ip1(n18296), .ip2(n18295), .op(n19320) );
  nand2_1 U22296 ( .ip1(n18297), .ip2(n19320), .op(n18302) );
  inv_1 U22297 ( .ip(n18298), .op(n18310) );
  nand2_1 U22298 ( .ip1(\x[42][13] ), .ip2(n24081), .op(n18300) );
  nand2_1 U22299 ( .ip1(\x[42][12] ), .ip2(n24233), .op(n18299) );
  nand2_1 U22300 ( .ip1(n18300), .ip2(n18299), .op(n18318) );
  nand2_1 U22301 ( .ip1(n18310), .ip2(n18318), .op(n18301) );
  nand4_1 U22302 ( .ip1(n18304), .ip2(n18303), .ip3(n18302), .ip4(n18301), 
        .op(n24869) );
  nand2_1 U22303 ( .ip1(n18306), .ip2(n18305), .op(n18307) );
  nand2_1 U22304 ( .ip1(n18308), .ip2(n18307), .op(n18332) );
  nor2_1 U22305 ( .ip1(n18310), .ip2(n18309), .op(n18323) );
  inv_1 U22306 ( .ip(n18311), .op(n18313) );
  nand2_1 U22307 ( .ip1(\x[42][8] ), .ip2(n24491), .op(n18312) );
  nand2_1 U22308 ( .ip1(n18313), .ip2(n18312), .op(n18315) );
  nand2_1 U22309 ( .ip1(n18315), .ip2(n18314), .op(n18317) );
  nand2_1 U22310 ( .ip1(n18317), .ip2(n18316), .op(n18320) );
  not_ab_or_c_or_d U22311 ( .ip1(n18321), .ip2(n18320), .ip3(n18319), .ip4(
        n18318), .op(n18322) );
  not_ab_or_c_or_d U22312 ( .ip1(n18325), .ip2(n18324), .ip3(n18323), .ip4(
        n18322), .op(n18331) );
  inv_1 U22313 ( .ip(n18326), .op(n18327) );
  nand3_1 U22314 ( .ip1(n18329), .ip2(n18328), .ip3(n18327), .op(n18330) );
  nand3_1 U22315 ( .ip1(n18332), .ip2(n18331), .ip3(n18330), .op(n24868) );
  nand2_1 U22316 ( .ip1(n24869), .ip2(n24868), .op(n24860) );
  nor2_1 U22317 ( .ip1(n24859), .ip2(n24860), .op(n24865) );
  or2_1 U22318 ( .ip1(n18334), .ip2(n18333), .op(n18337) );
  not_ab_or_c_or_d U22319 ( .ip1(n18338), .ip2(n18337), .ip3(n18336), .ip4(
        n18335), .op(n18356) );
  inv_1 U22320 ( .ip(n18339), .op(n18340) );
  nor2_1 U22321 ( .ip1(n18341), .ip2(n18340), .op(n18355) );
  inv_1 U22322 ( .ip(n18342), .op(n18345) );
  and2_1 U22323 ( .ip1(n18345), .ip2(n18343), .op(n18354) );
  nand2_1 U22324 ( .ip1(n18345), .ip2(n18344), .op(n18349) );
  or2_1 U22325 ( .ip1(n18346), .ip2(n18349), .op(n18352) );
  or2_1 U22326 ( .ip1(n18348), .ip2(n18347), .op(n18350) );
  or2_1 U22327 ( .ip1(n18350), .ip2(n18349), .op(n18351) );
  nand2_1 U22328 ( .ip1(n18352), .ip2(n18351), .op(n18353) );
  or4_1 U22329 ( .ip1(n18356), .ip2(n18355), .ip3(n18354), .ip4(n18353), .op(
        n24867) );
  nand2_1 U22330 ( .ip1(n24865), .ip2(n24867), .op(n24863) );
  nor2_1 U22331 ( .ip1(n24862), .ip2(n24863), .op(n24877) );
  or2_1 U22332 ( .ip1(n18358), .ip2(n18357), .op(n18377) );
  inv_1 U22333 ( .ip(n18359), .op(n18369) );
  inv_1 U22334 ( .ip(n18360), .op(n18362) );
  inv_1 U22335 ( .ip(n18361), .op(n18363) );
  or2_1 U22336 ( .ip1(n18362), .ip2(n18363), .op(n18366) );
  or2_1 U22337 ( .ip1(n18364), .ip2(n18363), .op(n18365) );
  nand2_1 U22338 ( .ip1(n18366), .ip2(n18365), .op(n18367) );
  not_ab_or_c_or_d U22339 ( .ip1(n18370), .ip2(n18369), .ip3(n18368), .ip4(
        n18367), .op(n18376) );
  inv_1 U22340 ( .ip(n18371), .op(n18373) );
  nand3_1 U22341 ( .ip1(n18374), .ip2(n18373), .ip3(n18372), .op(n18375) );
  nand3_1 U22342 ( .ip1(n18377), .ip2(n18376), .ip3(n18375), .op(n24878) );
  nand2_1 U22343 ( .ip1(n24877), .ip2(n24878), .op(n24875) );
  nor2_1 U22344 ( .ip1(n24874), .ip2(n24875), .op(n24887) );
  and2_1 U22345 ( .ip1(n24081), .ip2(\x[35][13] ), .op(n18378) );
  nor2_1 U22346 ( .ip1(\x[35][15] ), .ip2(n23143), .op(n18450) );
  not_ab_or_c_or_d U22347 ( .ip1(\x[35][14] ), .ip2(n24230), .ip3(n18378), 
        .ip4(n18450), .op(n18443) );
  nand2_1 U22348 ( .ip1(\x[35][12] ), .ip2(n24233), .op(n18379) );
  nand2_1 U22349 ( .ip1(n18443), .ip2(n18379), .op(n18436) );
  nand2_1 U22350 ( .ip1(\x[35][15] ), .ip2(n24186), .op(n18419) );
  nor2_1 U22351 ( .ip1(n17845), .ip2(n18380), .op(n18383) );
  nor4_1 U22352 ( .ip1(n18384), .ip2(n18383), .ip3(n18382), .ip4(n18381), .op(
        n18418) );
  nor2_1 U22353 ( .ip1(n24239), .ip2(\x[35][11] ), .op(n18386) );
  not_ab_or_c_or_d U22354 ( .ip1(\x[35][11] ), .ip2(n24456), .ip3(\x[35][10] ), 
        .ip4(n24370), .op(n18385) );
  or2_1 U22355 ( .ip1(n18386), .ip2(n18385), .op(n18432) );
  and2_1 U22356 ( .ip1(n24461), .ip2(\x[35][7] ), .op(n18402) );
  inv_1 U22357 ( .ip(\x[35][5] ), .op(n18400) );
  nor2_1 U22358 ( .ip1(n22833), .ip2(n18400), .op(n18397) );
  inv_1 U22359 ( .ip(\x[35][3] ), .op(n18395) );
  and2_1 U22360 ( .ip1(n24335), .ip2(\x[35][2] ), .op(n18392) );
  nand2_1 U22361 ( .ip1(\x[35][0] ), .ip2(n24143), .op(n18390) );
  nand2_1 U22362 ( .ip1(\x[35][1] ), .ip2(n20652), .op(n18389) );
  nor2_1 U22363 ( .ip1(\x[35][2] ), .ip2(n24463), .op(n18388) );
  nor2_1 U22364 ( .ip1(\x[35][1] ), .ip2(n21685), .op(n18387) );
  not_ab_or_c_or_d U22365 ( .ip1(n18390), .ip2(n18389), .ip3(n18388), .ip4(
        n18387), .op(n18391) );
  not_ab_or_c_or_d U22366 ( .ip1(\x[35][3] ), .ip2(n22795), .ip3(n18392), 
        .ip4(n18391), .op(n18394) );
  nor2_1 U22367 ( .ip1(\x[35][4] ), .ip2(n24256), .op(n18393) );
  not_ab_or_c_or_d U22368 ( .ip1(n23251), .ip2(n18395), .ip3(n18394), .ip4(
        n18393), .op(n18396) );
  not_ab_or_c_or_d U22369 ( .ip1(\x[35][4] ), .ip2(n23721), .ip3(n18397), 
        .ip4(n18396), .op(n18399) );
  nor2_1 U22370 ( .ip1(\x[35][6] ), .ip2(n23509), .op(n18398) );
  not_ab_or_c_or_d U22371 ( .ip1(sig_in[5]), .ip2(n18400), .ip3(n18399), .ip4(
        n18398), .op(n18401) );
  not_ab_or_c_or_d U22372 ( .ip1(\x[35][6] ), .ip2(n24355), .ip3(n18402), 
        .ip4(n18401), .op(n18404) );
  nor2_1 U22373 ( .ip1(\x[35][7] ), .ip2(n24142), .op(n18403) );
  nor2_1 U22374 ( .ip1(n18404), .ip2(n18403), .op(n18427) );
  buf_1 U22375 ( .ip(sig_in[8]), .op(n23779) );
  nor2_1 U22376 ( .ip1(\x[35][9] ), .ip2(n24043), .op(n18408) );
  or2_1 U22377 ( .ip1(n23779), .ip2(n18408), .op(n18407) );
  inv_1 U22378 ( .ip(\x[35][8] ), .op(n18405) );
  or2_1 U22379 ( .ip1(n18405), .ip2(n18408), .op(n18406) );
  nand2_1 U22380 ( .ip1(n18407), .ip2(n18406), .op(n18431) );
  nand2_1 U22381 ( .ip1(\x[35][8] ), .ip2(n23971), .op(n18428) );
  nor2_1 U22382 ( .ip1(n18408), .ip2(n18428), .op(n18412) );
  nand2_1 U22383 ( .ip1(n24455), .ip2(\x[35][9] ), .op(n18411) );
  nand2_1 U22384 ( .ip1(\x[35][11] ), .ip2(n21793), .op(n18410) );
  nand2_1 U22385 ( .ip1(\x[35][10] ), .ip2(n23980), .op(n18409) );
  nand3_1 U22386 ( .ip1(n18411), .ip2(n18410), .ip3(n18409), .op(n18425) );
  not_ab_or_c_or_d U22387 ( .ip1(n18427), .ip2(n18431), .ip3(n18412), .ip4(
        n18425), .op(n18416) );
  or2_1 U22388 ( .ip1(n24185), .ip2(\x[35][14] ), .op(n18413) );
  nand2_1 U22389 ( .ip1(n18419), .ip2(n18413), .op(n18448) );
  nor2_1 U22390 ( .ip1(\x[35][13] ), .ip2(n24332), .op(n18415) );
  nor2_1 U22391 ( .ip1(\x[35][12] ), .ip2(n24233), .op(n18414) );
  or2_1 U22392 ( .ip1(n18415), .ip2(n18414), .op(n18442) );
  nor4_1 U22393 ( .ip1(n18432), .ip2(n18416), .ip3(n18448), .ip4(n18442), .op(
        n18417) );
  not_ab_or_c_or_d U22394 ( .ip1(n18436), .ip2(n18419), .ip3(n18418), .ip4(
        n18417), .op(n18424) );
  inv_1 U22395 ( .ip(n18420), .op(n18421) );
  nand2_1 U22396 ( .ip1(n18422), .ip2(n18421), .op(n18423) );
  nand2_1 U22397 ( .ip1(n18424), .ip2(n18423), .op(n24892) );
  inv_1 U22398 ( .ip(n18425), .op(n18426) );
  or2_1 U22399 ( .ip1(n18426), .ip2(n18432), .op(n18435) );
  inv_1 U22400 ( .ip(n18427), .op(n18429) );
  nand2_1 U22401 ( .ip1(n18429), .ip2(n18428), .op(n18430) );
  nand2_1 U22402 ( .ip1(n18431), .ip2(n18430), .op(n18433) );
  or2_1 U22403 ( .ip1(n18433), .ip2(n18432), .op(n18434) );
  nand2_1 U22404 ( .ip1(n18435), .ip2(n18434), .op(n18437) );
  nor2_1 U22405 ( .ip1(n18437), .ip2(n18436), .op(n18441) );
  and2_1 U22406 ( .ip1(n18439), .ip2(n18438), .op(n18440) );
  not_ab_or_c_or_d U22407 ( .ip1(n18443), .ip2(n18442), .ip3(n18441), .ip4(
        n18440), .op(n18454) );
  nor2_1 U22408 ( .ip1(n18445), .ip2(n18444), .op(n18446) );
  nor2_1 U22409 ( .ip1(n18447), .ip2(n18446), .op(n18452) );
  inv_1 U22410 ( .ip(n18448), .op(n18449) );
  nor2_1 U22411 ( .ip1(n18450), .ip2(n18449), .op(n18451) );
  nor2_1 U22412 ( .ip1(n18452), .ip2(n18451), .op(n18453) );
  nand2_1 U22413 ( .ip1(n18454), .ip2(n18453), .op(n24888) );
  nand3_1 U22414 ( .ip1(n24887), .ip2(n24892), .ip3(n24888), .op(n24891) );
  nor3_1 U22415 ( .ip1(n24889), .ip2(n24880), .ip3(n24891), .op(n24853) );
  nor2_1 U22416 ( .ip1(n24384), .ip2(\x[31][15] ), .op(n18493) );
  nor2_1 U22417 ( .ip1(\x[31][12] ), .ip2(n24079), .op(n18485) );
  nor2_1 U22418 ( .ip1(\x[31][11] ), .ip2(n24239), .op(n18484) );
  nor2_1 U22419 ( .ip1(\x[31][13] ), .ip2(n24235), .op(n18483) );
  and2_1 U22420 ( .ip1(n24371), .ip2(\x[31][11] ), .op(n18479) );
  nor3_1 U22421 ( .ip1(n24370), .ip2(\x[31][10] ), .ip3(n18479), .op(n18481)
         );
  nor2_1 U22422 ( .ip1(\x[31][9] ), .ip2(n24043), .op(n18474) );
  inv_1 U22423 ( .ip(\x[31][8] ), .op(n18455) );
  nor3_1 U22424 ( .ip1(sig_in[8]), .ip2(n18474), .ip3(n18455), .op(n18477) );
  and2_1 U22425 ( .ip1(n24461), .ip2(\x[31][7] ), .op(n18471) );
  inv_1 U22426 ( .ip(\x[31][5] ), .op(n18469) );
  inv_1 U22427 ( .ip(n24462), .op(n23860) );
  nor2_1 U22428 ( .ip1(n22833), .ip2(n18469), .op(n18466) );
  inv_1 U22429 ( .ip(\x[31][3] ), .op(n18464) );
  and2_1 U22430 ( .ip1(n24335), .ip2(\x[31][2] ), .op(n18461) );
  nand2_1 U22431 ( .ip1(\x[31][1] ), .ip2(n21685), .op(n18459) );
  nand2_1 U22432 ( .ip1(\x[31][0] ), .ip2(n24143), .op(n18458) );
  nor2_1 U22433 ( .ip1(\x[31][2] ), .ip2(n24463), .op(n18457) );
  nor2_1 U22434 ( .ip1(\x[31][1] ), .ip2(n20652), .op(n18456) );
  not_ab_or_c_or_d U22435 ( .ip1(n18459), .ip2(n18458), .ip3(n18457), .ip4(
        n18456), .op(n18460) );
  not_ab_or_c_or_d U22436 ( .ip1(\x[31][3] ), .ip2(n22795), .ip3(n18461), 
        .ip4(n18460), .op(n18463) );
  nor2_1 U22437 ( .ip1(\x[31][4] ), .ip2(n24256), .op(n18462) );
  not_ab_or_c_or_d U22438 ( .ip1(n23251), .ip2(n18464), .ip3(n18463), .ip4(
        n18462), .op(n18465) );
  not_ab_or_c_or_d U22439 ( .ip1(\x[31][4] ), .ip2(n23860), .ip3(n18466), 
        .ip4(n18465), .op(n18468) );
  nor2_1 U22440 ( .ip1(\x[31][6] ), .ip2(n23770), .op(n18467) );
  not_ab_or_c_or_d U22441 ( .ip1(sig_in[5]), .ip2(n18469), .ip3(n18468), .ip4(
        n18467), .op(n18470) );
  not_ab_or_c_or_d U22442 ( .ip1(\x[31][6] ), .ip2(n24355), .ip3(n18471), 
        .ip4(n18470), .op(n18475) );
  nor2_1 U22443 ( .ip1(\x[31][8] ), .ip2(n24358), .op(n18473) );
  nor2_1 U22444 ( .ip1(\x[31][7] ), .ip2(n24492), .op(n18472) );
  nor4_1 U22445 ( .ip1(n18475), .ip2(n18474), .ip3(n18473), .ip4(n18472), .op(
        n18476) );
  ab_or_c_or_d U22446 ( .ip1(\x[31][9] ), .ip2(n24043), .ip3(n18477), .ip4(
        n18476), .op(n18478) );
  not_ab_or_c_or_d U22447 ( .ip1(\x[31][10] ), .ip2(n20880), .ip3(n18479), 
        .ip4(n18478), .op(n18480) );
  or2_1 U22448 ( .ip1(n18481), .ip2(n18480), .op(n18482) );
  nor4_1 U22449 ( .ip1(n18485), .ip2(n18484), .ip3(n18483), .ip4(n18482), .op(
        n18489) );
  nand2_1 U22450 ( .ip1(\x[31][13] ), .ip2(n24235), .op(n18487) );
  nand2_1 U22451 ( .ip1(\x[31][12] ), .ip2(n24449), .op(n18486) );
  nand2_1 U22452 ( .ip1(n18487), .ip2(n18486), .op(n18488) );
  not_ab_or_c_or_d U22453 ( .ip1(\x[31][14] ), .ip2(n24230), .ip3(n18489), 
        .ip4(n18488), .op(n18491) );
  nor2_1 U22454 ( .ip1(\x[31][14] ), .ip2(n23938), .op(n18490) );
  not_ab_or_c_or_d U22455 ( .ip1(\x[31][15] ), .ip2(n24384), .ip3(n18491), 
        .ip4(n18490), .op(n18492) );
  or2_1 U22456 ( .ip1(n18493), .ip2(n18492), .op(n18503) );
  nand2_1 U22457 ( .ip1(n18494), .ip2(n18503), .op(n24855) );
  or2_1 U22458 ( .ip1(n18495), .ip2(n18498), .op(n18501) );
  nand2_1 U22459 ( .ip1(n18497), .ip2(n18496), .op(n18499) );
  or2_1 U22460 ( .ip1(n18499), .ip2(n18498), .op(n18500) );
  nand2_1 U22461 ( .ip1(n18501), .ip2(n18500), .op(n18502) );
  ab_or_c_or_d U22462 ( .ip1(n18505), .ip2(n18504), .ip3(n18503), .ip4(n18502), 
        .op(n24854) );
  nand3_1 U22463 ( .ip1(n24853), .ip2(n24855), .ip3(n24854), .op(n24852) );
  nor2_1 U22464 ( .ip1(\x[58][15] ), .ip2(n23143), .op(n18554) );
  or2_1 U22465 ( .ip1(\x[58][14] ), .ip2(n18554), .op(n18507) );
  or2_1 U22466 ( .ip1(n24230), .ip2(n18554), .op(n18506) );
  nand2_1 U22467 ( .ip1(n18507), .ip2(n18506), .op(n18599) );
  inv_1 U22468 ( .ip(\x[58][12] ), .op(n18550) );
  and2_1 U22469 ( .ip1(n24235), .ip2(\x[58][13] ), .op(n18547) );
  nand2_1 U22470 ( .ip1(\x[58][10] ), .ip2(n23980), .op(n18537) );
  inv_1 U22471 ( .ip(n21171), .op(n23981) );
  nor2_1 U22472 ( .ip1(\x[58][9] ), .ip2(n24455), .op(n18532) );
  inv_1 U22473 ( .ip(\x[58][8] ), .op(n18508) );
  nor3_1 U22474 ( .ip1(sig_in[8]), .ip2(n18532), .ip3(n18508), .op(n18535) );
  and2_1 U22475 ( .ip1(n24461), .ip2(\x[58][7] ), .op(n18529) );
  inv_1 U22476 ( .ip(\x[58][5] ), .op(n18527) );
  nor2_1 U22477 ( .ip1(n22833), .ip2(n18527), .op(n18524) );
  inv_1 U22478 ( .ip(\x[58][3] ), .op(n18515) );
  inv_1 U22479 ( .ip(\x[58][1] ), .op(n18510) );
  nor2_1 U22480 ( .ip1(n24467), .ip2(n18510), .op(n18512) );
  inv_1 U22481 ( .ip(\x[58][0] ), .op(n18509) );
  not_ab_or_c_or_d U22482 ( .ip1(n22513), .ip2(n18510), .ip3(sig_in[0]), .ip4(
        n18509), .op(n18511) );
  not_ab_or_c_or_d U22483 ( .ip1(\x[58][2] ), .ip2(n24335), .ip3(n18512), 
        .ip4(n18511), .op(n18514) );
  nor2_1 U22484 ( .ip1(\x[58][2] ), .ip2(n24463), .op(n18513) );
  not_ab_or_c_or_d U22485 ( .ip1(n24251), .ip2(n18515), .ip3(n18514), .ip4(
        n18513), .op(n18516) );
  or2_1 U22486 ( .ip1(\x[58][3] ), .ip2(n18516), .op(n18518) );
  or2_1 U22487 ( .ip1(n22795), .ip2(n18516), .op(n18517) );
  nand2_1 U22488 ( .ip1(n18518), .ip2(n18517), .op(n18519) );
  or2_1 U22489 ( .ip1(sig_in[4]), .ip2(n18519), .op(n18522) );
  inv_1 U22490 ( .ip(\x[58][4] ), .op(n18520) );
  or2_1 U22491 ( .ip1(n18520), .ip2(n18519), .op(n18521) );
  nand2_1 U22492 ( .ip1(n18522), .ip2(n18521), .op(n18523) );
  not_ab_or_c_or_d U22493 ( .ip1(\x[58][4] ), .ip2(n23860), .ip3(n18524), 
        .ip4(n18523), .op(n18526) );
  nor2_1 U22494 ( .ip1(\x[58][6] ), .ip2(n23770), .op(n18525) );
  not_ab_or_c_or_d U22495 ( .ip1(sig_in[5]), .ip2(n18527), .ip3(n18526), .ip4(
        n18525), .op(n18528) );
  not_ab_or_c_or_d U22496 ( .ip1(\x[58][6] ), .ip2(n24485), .ip3(n18529), 
        .ip4(n18528), .op(n18533) );
  nor2_1 U22497 ( .ip1(\x[58][7] ), .ip2(n24492), .op(n18531) );
  nor2_1 U22498 ( .ip1(\x[58][8] ), .ip2(n24358), .op(n18530) );
  nor4_1 U22499 ( .ip1(n18533), .ip2(n18532), .ip3(n18531), .ip4(n18530), .op(
        n18534) );
  not_ab_or_c_or_d U22500 ( .ip1(\x[58][9] ), .ip2(n23981), .ip3(n18535), 
        .ip4(n18534), .op(n18536) );
  nand2_1 U22501 ( .ip1(n18537), .ip2(n18536), .op(n18543) );
  nor2_1 U22502 ( .ip1(\x[58][10] ), .ip2(n20880), .op(n18538) );
  or2_1 U22503 ( .ip1(sig_in[11]), .ip2(n18538), .op(n18541) );
  inv_1 U22504 ( .ip(\x[58][11] ), .op(n18539) );
  or2_1 U22505 ( .ip1(n18539), .ip2(n18538), .op(n18540) );
  nand2_1 U22506 ( .ip1(n18541), .ip2(n18540), .op(n18542) );
  nand2_1 U22507 ( .ip1(n18543), .ip2(n18542), .op(n18545) );
  nand2_1 U22508 ( .ip1(\x[58][11] ), .ip2(n24456), .op(n18544) );
  nand2_1 U22509 ( .ip1(n18545), .ip2(n18544), .op(n18546) );
  not_ab_or_c_or_d U22510 ( .ip1(\x[58][12] ), .ip2(n24079), .ip3(n18547), 
        .ip4(n18546), .op(n18549) );
  nor2_1 U22511 ( .ip1(\x[58][13] ), .ip2(n24137), .op(n18548) );
  not_ab_or_c_or_d U22512 ( .ip1(n17845), .ip2(n18550), .ip3(n18549), .ip4(
        n18548), .op(n18653) );
  inv_1 U22513 ( .ip(n18653), .op(n18598) );
  and2_1 U22514 ( .ip1(n24186), .ip2(\x[58][15] ), .op(n18600) );
  or2_1 U22515 ( .ip1(sig_in[14]), .ip2(n18600), .op(n18553) );
  inv_1 U22516 ( .ip(\x[58][14] ), .op(n18551) );
  or2_1 U22517 ( .ip1(n18551), .ip2(n18600), .op(n18552) );
  nand2_1 U22518 ( .ip1(n18553), .ip2(n18552), .op(n18652) );
  nor2_1 U22519 ( .ip1(n18652), .ip2(n18554), .op(n18597) );
  nor2_1 U22520 ( .ip1(n24384), .ip2(\x[57][15] ), .op(n18596) );
  and2_1 U22521 ( .ip1(n24081), .ip2(\x[57][13] ), .op(n18587) );
  and2_1 U22522 ( .ip1(n24461), .ip2(\x[57][7] ), .op(n18571) );
  inv_1 U22523 ( .ip(\x[57][3] ), .op(n18561) );
  inv_1 U22524 ( .ip(\x[57][1] ), .op(n18556) );
  nor2_1 U22525 ( .ip1(n22513), .ip2(n18556), .op(n18558) );
  inv_1 U22526 ( .ip(\x[57][0] ), .op(n18555) );
  not_ab_or_c_or_d U22527 ( .ip1(n22513), .ip2(n18556), .ip3(sig_in[0]), .ip4(
        n18555), .op(n18557) );
  not_ab_or_c_or_d U22528 ( .ip1(\x[57][2] ), .ip2(n24470), .ip3(n18558), 
        .ip4(n18557), .op(n18560) );
  nor2_1 U22529 ( .ip1(\x[57][2] ), .ip2(n24463), .op(n18559) );
  not_ab_or_c_or_d U22530 ( .ip1(n23251), .ip2(n18561), .ip3(n18560), .ip4(
        n18559), .op(n18565) );
  buf_1 U22531 ( .ip(n23283), .op(n24119) );
  nand2_1 U22532 ( .ip1(\x[57][5] ), .ip2(n24119), .op(n18563) );
  nand2_1 U22533 ( .ip1(\x[57][4] ), .ip2(n23721), .op(n18562) );
  nand2_1 U22534 ( .ip1(n18563), .ip2(n18562), .op(n18564) );
  not_ab_or_c_or_d U22535 ( .ip1(\x[57][3] ), .ip2(n22795), .ip3(n18565), 
        .ip4(n18564), .op(n18569) );
  nor2_1 U22536 ( .ip1(\x[57][5] ), .ip2(n23283), .op(n18568) );
  nor2_1 U22537 ( .ip1(\x[57][6] ), .ip2(n24355), .op(n18567) );
  not_ab_or_c_or_d U22538 ( .ip1(\x[57][5] ), .ip2(n23600), .ip3(\x[57][4] ), 
        .ip4(n24347), .op(n18566) );
  nor4_1 U22539 ( .ip1(n18569), .ip2(n18568), .ip3(n18567), .ip4(n18566), .op(
        n18570) );
  not_ab_or_c_or_d U22540 ( .ip1(\x[57][6] ), .ip2(n23770), .ip3(n18571), 
        .ip4(n18570), .op(n18574) );
  nor2_1 U22541 ( .ip1(\x[57][9] ), .ip2(n24455), .op(n18575) );
  nor2_1 U22542 ( .ip1(\x[57][8] ), .ip2(n23971), .op(n18573) );
  nor2_1 U22543 ( .ip1(\x[57][7] ), .ip2(n24142), .op(n18572) );
  nor4_1 U22544 ( .ip1(n18574), .ip2(n18575), .ip3(n18573), .ip4(n18572), .op(
        n18581) );
  nand2_1 U22545 ( .ip1(n24455), .ip2(\x[57][9] ), .op(n18579) );
  inv_1 U22546 ( .ip(n18575), .op(n18576) );
  nand3_1 U22547 ( .ip1(\x[57][8] ), .ip2(n24100), .ip3(n18576), .op(n18578)
         );
  nand2_1 U22548 ( .ip1(\x[57][11] ), .ip2(n24456), .op(n18577) );
  nand3_1 U22549 ( .ip1(n18579), .ip2(n18578), .ip3(n18577), .op(n18580) );
  not_ab_or_c_or_d U22550 ( .ip1(\x[57][10] ), .ip2(n23980), .ip3(n18581), 
        .ip4(n18580), .op(n18585) );
  nor2_1 U22551 ( .ip1(\x[57][11] ), .ip2(n24371), .op(n18584) );
  nor2_1 U22552 ( .ip1(\x[57][12] ), .ip2(n24233), .op(n18583) );
  not_ab_or_c_or_d U22553 ( .ip1(\x[57][11] ), .ip2(n24136), .ip3(\x[57][10] ), 
        .ip4(n20880), .op(n18582) );
  nor4_1 U22554 ( .ip1(n18585), .ip2(n18584), .ip3(n18583), .ip4(n18582), .op(
        n18586) );
  not_ab_or_c_or_d U22555 ( .ip1(\x[57][12] ), .ip2(n24079), .ip3(n18587), 
        .ip4(n18586), .op(n18589) );
  nor2_1 U22556 ( .ip1(\x[57][13] ), .ip2(n24376), .op(n18588) );
  nor2_1 U22557 ( .ip1(n18589), .ip2(n18588), .op(n18590) );
  or2_1 U22558 ( .ip1(\x[57][14] ), .ip2(n18590), .op(n18592) );
  or2_1 U22559 ( .ip1(n24230), .ip2(n18590), .op(n18591) );
  nand2_1 U22560 ( .ip1(n18592), .ip2(n18591), .op(n18594) );
  nor2_1 U22561 ( .ip1(\x[57][14] ), .ip2(n23938), .op(n18593) );
  not_ab_or_c_or_d U22562 ( .ip1(\x[57][15] ), .ip2(n24384), .ip3(n18594), 
        .ip4(n18593), .op(n18595) );
  or2_1 U22563 ( .ip1(n18596), .ip2(n18595), .op(n19941) );
  not_ab_or_c_or_d U22564 ( .ip1(n18599), .ip2(n18598), .ip3(n18597), .ip4(
        n19941), .op(n24683) );
  nor2_1 U22565 ( .ip1(n18600), .ip2(n18599), .op(n18651) );
  nor2_1 U22566 ( .ip1(\x[59][14] ), .ip2(n23938), .op(n18601) );
  or2_1 U22567 ( .ip1(\x[59][15] ), .ip2(n18601), .op(n18603) );
  or2_1 U22568 ( .ip1(n24329), .ip2(n18601), .op(n18602) );
  nand2_1 U22569 ( .ip1(n18603), .ip2(n18602), .op(n18650) );
  nand2_1 U22570 ( .ip1(\x[59][13] ), .ip2(n24081), .op(n18605) );
  nand2_1 U22571 ( .ip1(\x[59][14] ), .ip2(n24327), .op(n18604) );
  nand2_1 U22572 ( .ip1(n18605), .ip2(n18604), .op(n18649) );
  nor2_1 U22573 ( .ip1(\x[59][15] ), .ip2(n23143), .op(n18648) );
  inv_1 U22574 ( .ip(\x[59][9] ), .op(n18626) );
  nand2_1 U22575 ( .ip1(n21171), .ip2(n18626), .op(n18632) );
  inv_1 U22576 ( .ip(\x[59][10] ), .op(n18633) );
  not_ab_or_c_or_d U22577 ( .ip1(\x[59][9] ), .ip2(n24043), .ip3(\x[59][8] ), 
        .ip4(n24358), .op(n18630) );
  and2_1 U22578 ( .ip1(n24461), .ip2(\x[59][7] ), .op(n18623) );
  nor2_1 U22579 ( .ip1(n23509), .ip2(\x[59][6] ), .op(n18621) );
  and2_1 U22580 ( .ip1(n23283), .ip2(\x[59][5] ), .op(n18619) );
  nor2_1 U22581 ( .ip1(\x[59][4] ), .ip2(n24347), .op(n18617) );
  and2_1 U22582 ( .ip1(n24347), .ip2(\x[59][4] ), .op(n18614) );
  inv_1 U22583 ( .ip(\x[59][3] ), .op(n18612) );
  nor2_1 U22584 ( .ip1(\x[59][2] ), .ip2(n24463), .op(n18611) );
  inv_1 U22585 ( .ip(\x[59][1] ), .op(n18607) );
  nor2_1 U22586 ( .ip1(n22513), .ip2(n18607), .op(n18609) );
  inv_1 U22587 ( .ip(\x[59][0] ), .op(n18606) );
  not_ab_or_c_or_d U22588 ( .ip1(n22513), .ip2(n18607), .ip3(sig_in[0]), .ip4(
        n18606), .op(n18608) );
  not_ab_or_c_or_d U22589 ( .ip1(\x[59][2] ), .ip2(n24335), .ip3(n18609), 
        .ip4(n18608), .op(n18610) );
  not_ab_or_c_or_d U22590 ( .ip1(n24251), .ip2(n18612), .ip3(n18611), .ip4(
        n18610), .op(n18613) );
  not_ab_or_c_or_d U22591 ( .ip1(\x[59][3] ), .ip2(n22795), .ip3(n18614), 
        .ip4(n18613), .op(n18616) );
  nor2_1 U22592 ( .ip1(\x[59][5] ), .ip2(n24119), .op(n18615) );
  nor3_1 U22593 ( .ip1(n18617), .ip2(n18616), .ip3(n18615), .op(n18618) );
  nor2_1 U22594 ( .ip1(n18619), .ip2(n18618), .op(n18620) );
  nor2_1 U22595 ( .ip1(n18621), .ip2(n18620), .op(n18622) );
  not_ab_or_c_or_d U22596 ( .ip1(\x[59][6] ), .ip2(n23509), .ip3(n18623), 
        .ip4(n18622), .op(n18625) );
  nor2_1 U22597 ( .ip1(\x[59][7] ), .ip2(n24044), .op(n18624) );
  nor2_1 U22598 ( .ip1(n18625), .ip2(n18624), .op(n18628) );
  nor2_1 U22599 ( .ip1(n21171), .ip2(n18626), .op(n18627) );
  not_ab_or_c_or_d U22600 ( .ip1(\x[59][8] ), .ip2(n24491), .ip3(n18628), 
        .ip4(n18627), .op(n18629) );
  not_ab_or_c_or_d U22601 ( .ip1(sig_in[10]), .ip2(n18633), .ip3(n18630), 
        .ip4(n18629), .op(n18631) );
  nand2_1 U22602 ( .ip1(n18632), .ip2(n18631), .op(n18638) );
  nor2_1 U22603 ( .ip1(sig_in[10]), .ip2(n18633), .op(n18634) );
  or2_1 U22604 ( .ip1(\x[59][11] ), .ip2(n18634), .op(n18636) );
  or2_1 U22605 ( .ip1(n24136), .ip2(n18634), .op(n18635) );
  nand2_1 U22606 ( .ip1(n18636), .ip2(n18635), .op(n18637) );
  nand2_1 U22607 ( .ip1(n18638), .ip2(n18637), .op(n18640) );
  or2_1 U22608 ( .ip1(n24239), .ip2(\x[59][11] ), .op(n18639) );
  nand2_1 U22609 ( .ip1(n18640), .ip2(n18639), .op(n18644) );
  or2_1 U22610 ( .ip1(n24081), .ip2(\x[59][13] ), .op(n18641) );
  nand2_1 U22611 ( .ip1(n18650), .ip2(n18641), .op(n18642) );
  nor3_1 U22612 ( .ip1(n18644), .ip2(n17845), .ip3(n18642), .op(n18646) );
  inv_1 U22613 ( .ip(\x[59][12] ), .op(n18643) );
  not_ab_or_c_or_d U22614 ( .ip1(n18644), .ip2(n17845), .ip3(n18643), .ip4(
        n18642), .op(n18645) );
  or2_1 U22615 ( .ip1(n18646), .ip2(n18645), .op(n18647) );
  not_ab_or_c_or_d U22616 ( .ip1(n18650), .ip2(n18649), .ip3(n18648), .ip4(
        n18647), .op(n19316) );
  not_ab_or_c_or_d U22617 ( .ip1(n18653), .ip2(n18652), .ip3(n18651), .ip4(
        n19316), .op(n24651) );
  and2_1 U22618 ( .ip1(n23895), .ip2(\x[60][13] ), .op(n18654) );
  nor2_1 U22619 ( .ip1(\x[60][15] ), .ip2(n23143), .op(n19307) );
  not_ab_or_c_or_d U22620 ( .ip1(\x[60][14] ), .ip2(n24230), .ip3(n18654), 
        .ip4(n19307), .op(n19314) );
  nand2_1 U22621 ( .ip1(\x[60][12] ), .ip2(n24450), .op(n19311) );
  nand2_1 U22622 ( .ip1(n19314), .ip2(n19311), .op(n18749) );
  nand2_1 U22623 ( .ip1(\x[60][15] ), .ip2(n24186), .op(n18748) );
  nor2_1 U22624 ( .ip1(\x[61][11] ), .ip2(n21793), .op(n19279) );
  nor2_1 U22625 ( .ip1(\x[61][10] ), .ip2(n20880), .op(n18655) );
  nor2_1 U22626 ( .ip1(n19279), .ip2(n18655), .op(n19288) );
  inv_1 U22627 ( .ip(n19288), .op(n19280) );
  nor2_1 U22628 ( .ip1(\x[61][9] ), .ip2(n24269), .op(n19281) );
  or2_1 U22629 ( .ip1(n23779), .ip2(n19281), .op(n18658) );
  inv_1 U22630 ( .ip(\x[61][8] ), .op(n18656) );
  or2_1 U22631 ( .ip1(n18656), .ip2(n19281), .op(n18657) );
  nand2_1 U22632 ( .ip1(n18658), .ip2(n18657), .op(n19289) );
  nor2_1 U22633 ( .ip1(n24142), .ip2(\x[61][7] ), .op(n18681) );
  inv_1 U22634 ( .ip(\x[61][5] ), .op(n18677) );
  inv_1 U22635 ( .ip(\x[61][4] ), .op(n18669) );
  nor2_1 U22636 ( .ip1(n24462), .ip2(n18669), .op(n18667) );
  inv_1 U22637 ( .ip(\x[61][3] ), .op(n18665) );
  inv_1 U22638 ( .ip(\x[61][1] ), .op(n18660) );
  nor2_1 U22639 ( .ip1(n22513), .ip2(n18660), .op(n18662) );
  inv_1 U22640 ( .ip(\x[61][0] ), .op(n18659) );
  not_ab_or_c_or_d U22641 ( .ip1(n24467), .ip2(n18660), .ip3(sig_in[0]), .ip4(
        n18659), .op(n18661) );
  not_ab_or_c_or_d U22642 ( .ip1(\x[61][2] ), .ip2(n24470), .ip3(n18662), 
        .ip4(n18661), .op(n18664) );
  nor2_1 U22643 ( .ip1(\x[61][2] ), .ip2(n24463), .op(n18663) );
  not_ab_or_c_or_d U22644 ( .ip1(n24251), .ip2(n18665), .ip3(n18664), .ip4(
        n18663), .op(n18666) );
  not_ab_or_c_or_d U22645 ( .ip1(\x[61][3] ), .ip2(n22795), .ip3(n18667), 
        .ip4(n18666), .op(n18668) );
  or2_1 U22646 ( .ip1(sig_in[4]), .ip2(n18668), .op(n18671) );
  or2_1 U22647 ( .ip1(n18669), .ip2(n18668), .op(n18670) );
  nand2_1 U22648 ( .ip1(n18671), .ip2(n18670), .op(n18672) );
  or2_1 U22649 ( .ip1(\x[61][5] ), .ip2(n18672), .op(n18674) );
  or2_1 U22650 ( .ip1(n23600), .ip2(n18672), .op(n18673) );
  nand2_1 U22651 ( .ip1(n18674), .ip2(n18673), .op(n18676) );
  nor2_1 U22652 ( .ip1(\x[61][6] ), .ip2(n23509), .op(n18675) );
  not_ab_or_c_or_d U22653 ( .ip1(n22833), .ip2(n18677), .ip3(n18676), .ip4(
        n18675), .op(n18679) );
  and2_1 U22654 ( .ip1(n23770), .ip2(\x[61][6] ), .op(n18678) );
  not_ab_or_c_or_d U22655 ( .ip1(\x[61][7] ), .ip2(n24044), .ip3(n18679), 
        .ip4(n18678), .op(n18680) );
  nor2_1 U22656 ( .ip1(n18681), .ip2(n18680), .op(n19290) );
  inv_1 U22657 ( .ip(n19290), .op(n18682) );
  nand2_1 U22658 ( .ip1(\x[61][8] ), .ip2(n23804), .op(n19283) );
  nand2_1 U22659 ( .ip1(n18682), .ip2(n19283), .op(n18685) );
  nand2_1 U22660 ( .ip1(n24455), .ip2(\x[61][9] ), .op(n19282) );
  inv_1 U22661 ( .ip(n19282), .op(n18684) );
  nand2_1 U22662 ( .ip1(\x[61][11] ), .ip2(n21793), .op(n18687) );
  nand2_1 U22663 ( .ip1(\x[61][10] ), .ip2(n23980), .op(n18683) );
  nand2_1 U22664 ( .ip1(n18687), .ip2(n18683), .op(n19286) );
  not_ab_or_c_or_d U22665 ( .ip1(n19289), .ip2(n18685), .ip3(n18684), .ip4(
        n19286), .op(n18686) );
  or2_1 U22666 ( .ip1(n19280), .ip2(n18686), .op(n18688) );
  nand2_1 U22667 ( .ip1(n18688), .ip2(n18687), .op(n18692) );
  and2_1 U22668 ( .ip1(n24332), .ip2(\x[61][13] ), .op(n18690) );
  nor2_1 U22669 ( .ip1(\x[61][15] ), .ip2(n23143), .op(n18689) );
  not_ab_or_c_or_d U22670 ( .ip1(\x[61][14] ), .ip2(n24185), .ip3(n18690), 
        .ip4(n18689), .op(n18696) );
  nand2_1 U22671 ( .ip1(\x[61][12] ), .ip2(n24079), .op(n18691) );
  nand2_1 U22672 ( .ip1(n18696), .ip2(n18691), .op(n19284) );
  nor2_1 U22673 ( .ip1(n18692), .ip2(n19284), .op(n18747) );
  inv_1 U22674 ( .ip(\x[61][15] ), .op(n18693) );
  nor2_1 U22675 ( .ip1(n18693), .ip2(sig_in[15]), .op(n18695) );
  not_ab_or_c_or_d U22676 ( .ip1(sig_in[15]), .ip2(n18693), .ip3(\x[61][14] ), 
        .ip4(n24230), .op(n18694) );
  or2_1 U22677 ( .ip1(n18695), .ip2(n18694), .op(n18699) );
  or2_1 U22678 ( .ip1(n18696), .ip2(n18699), .op(n18702) );
  nor2_1 U22679 ( .ip1(\x[61][13] ), .ip2(n24081), .op(n18698) );
  nor2_1 U22680 ( .ip1(\x[61][12] ), .ip2(n24233), .op(n18697) );
  or2_1 U22681 ( .ip1(n18698), .ip2(n18697), .op(n18700) );
  or2_1 U22682 ( .ip1(n18700), .ip2(n18699), .op(n18701) );
  nand2_1 U22683 ( .ip1(n18702), .ip2(n18701), .op(n19294) );
  nor2_1 U22684 ( .ip1(\x[60][13] ), .ip2(n23895), .op(n18703) );
  or2_1 U22685 ( .ip1(n17845), .ip2(n18703), .op(n18706) );
  inv_1 U22686 ( .ip(\x[60][12] ), .op(n18704) );
  or2_1 U22687 ( .ip1(n18704), .ip2(n18703), .op(n18705) );
  nand2_1 U22688 ( .ip1(n18706), .ip2(n18705), .op(n19312) );
  inv_1 U22689 ( .ip(n18748), .op(n18707) );
  or2_1 U22690 ( .ip1(sig_in[14]), .ip2(n18707), .op(n18710) );
  inv_1 U22691 ( .ip(\x[60][14] ), .op(n18708) );
  or2_1 U22692 ( .ip1(n18708), .ip2(n18707), .op(n18709) );
  nand2_1 U22693 ( .ip1(n18710), .ip2(n18709), .op(n19308) );
  and2_1 U22694 ( .ip1(n24371), .ip2(\x[60][11] ), .op(n18737) );
  and2_1 U22695 ( .ip1(n24335), .ip2(\x[60][2] ), .op(n18716) );
  nand2_1 U22696 ( .ip1(\x[60][1] ), .ip2(n20652), .op(n18714) );
  nand2_1 U22697 ( .ip1(\x[60][0] ), .ip2(n24143), .op(n18713) );
  nor2_1 U22698 ( .ip1(\x[60][2] ), .ip2(n24463), .op(n18712) );
  nor2_1 U22699 ( .ip1(\x[60][1] ), .ip2(n21685), .op(n18711) );
  not_ab_or_c_or_d U22700 ( .ip1(n18714), .ip2(n18713), .ip3(n18712), .ip4(
        n18711), .op(n18715) );
  not_ab_or_c_or_d U22701 ( .ip1(\x[60][3] ), .ip2(n22795), .ip3(n18716), 
        .ip4(n18715), .op(n18719) );
  nor2_1 U22702 ( .ip1(\x[60][5] ), .ip2(n23283), .op(n18720) );
  nor2_1 U22703 ( .ip1(\x[60][4] ), .ip2(n23860), .op(n18718) );
  nor2_1 U22704 ( .ip1(\x[60][3] ), .ip2(n24342), .op(n18717) );
  nor4_1 U22705 ( .ip1(n18719), .ip2(n18720), .ip3(n18718), .ip4(n18717), .op(
        n18726) );
  nand2_1 U22706 ( .ip1(n23600), .ip2(\x[60][5] ), .op(n18724) );
  inv_1 U22707 ( .ip(n18720), .op(n18721) );
  nand3_1 U22708 ( .ip1(\x[60][4] ), .ip2(n23721), .ip3(n18721), .op(n18723)
         );
  inv_1 U22709 ( .ip(n17732), .op(n24044) );
  nand2_1 U22710 ( .ip1(\x[60][7] ), .ip2(n24044), .op(n18722) );
  nand3_1 U22711 ( .ip1(n18724), .ip2(n18723), .ip3(n18722), .op(n18725) );
  not_ab_or_c_or_d U22712 ( .ip1(\x[60][6] ), .ip2(n24355), .ip3(n18726), 
        .ip4(n18725), .op(n18730) );
  not_ab_or_c_or_d U22713 ( .ip1(\x[60][7] ), .ip2(n24142), .ip3(\x[60][6] ), 
        .ip4(n23770), .op(n18729) );
  nor2_1 U22714 ( .ip1(\x[60][7] ), .ip2(n24142), .op(n18728) );
  nor2_1 U22715 ( .ip1(\x[60][8] ), .ip2(n23971), .op(n18727) );
  or4_1 U22716 ( .ip1(n18730), .ip2(n18729), .ip3(n18728), .ip4(n18727), .op(
        n18731) );
  nor2_1 U22717 ( .ip1(\x[60][9] ), .ip2(n24164), .op(n18732) );
  or2_1 U22718 ( .ip1(n18731), .ip2(n18732), .op(n18735) );
  nand2_1 U22719 ( .ip1(\x[60][8] ), .ip2(n24100), .op(n18733) );
  or2_1 U22720 ( .ip1(n18733), .ip2(n18732), .op(n18734) );
  nand2_1 U22721 ( .ip1(n18735), .ip2(n18734), .op(n18736) );
  not_ab_or_c_or_d U22722 ( .ip1(\x[60][10] ), .ip2(n20880), .ip3(n18737), 
        .ip4(n18736), .op(n18740) );
  nor2_1 U22723 ( .ip1(n21793), .ip2(\x[60][11] ), .op(n18739) );
  not_ab_or_c_or_d U22724 ( .ip1(\x[60][11] ), .ip2(n24136), .ip3(\x[60][10] ), 
        .ip4(n24370), .op(n18738) );
  or2_1 U22725 ( .ip1(n18739), .ip2(n18738), .op(n18741) );
  or2_1 U22726 ( .ip1(n18740), .ip2(n18741), .op(n18744) );
  nand2_1 U22727 ( .ip1(\x[60][9] ), .ip2(n24043), .op(n18742) );
  or2_1 U22728 ( .ip1(n18742), .ip2(n18741), .op(n18743) );
  nand2_1 U22729 ( .ip1(n18744), .ip2(n18743), .op(n19309) );
  nand3_1 U22730 ( .ip1(n19312), .ip2(n19308), .ip3(n19309), .op(n18745) );
  nand2_1 U22731 ( .ip1(n19294), .ip2(n18745), .op(n18746) );
  not_ab_or_c_or_d U22732 ( .ip1(n18749), .ip2(n18748), .ip3(n18747), .ip4(
        n18746), .op(n24691) );
  and2_1 U22733 ( .ip1(n23895), .ip2(\x[66][13] ), .op(n18750) );
  nor2_1 U22734 ( .ip1(\x[66][15] ), .ip2(n23143), .op(n18756) );
  not_ab_or_c_or_d U22735 ( .ip1(\x[66][14] ), .ip2(n24185), .ip3(n18750), 
        .ip4(n18756), .op(n18841) );
  nor2_1 U22736 ( .ip1(\x[66][13] ), .ip2(n24332), .op(n18752) );
  nor2_1 U22737 ( .ip1(\x[66][12] ), .ip2(n24079), .op(n18751) );
  nor2_1 U22738 ( .ip1(n18752), .ip2(n18751), .op(n19114) );
  inv_1 U22739 ( .ip(n19114), .op(n18840) );
  nor2_1 U22740 ( .ip1(\x[66][14] ), .ip2(n23938), .op(n18753) );
  or2_1 U22741 ( .ip1(\x[66][15] ), .ip2(n18753), .op(n18755) );
  or2_1 U22742 ( .ip1(n24384), .ip2(n18753), .op(n18754) );
  nand2_1 U22743 ( .ip1(n18755), .ip2(n18754), .op(n19115) );
  nor2_1 U22744 ( .ip1(n18756), .ip2(n19115), .op(n19104) );
  and2_1 U22745 ( .ip1(n24332), .ip2(\x[65][13] ), .op(n18757) );
  nor2_1 U22746 ( .ip1(\x[65][15] ), .ip2(n23143), .op(n19173) );
  not_ab_or_c_or_d U22747 ( .ip1(\x[65][14] ), .ip2(n24185), .ip3(n18757), 
        .ip4(n19173), .op(n19168) );
  nand2_1 U22748 ( .ip1(\x[65][12] ), .ip2(n24233), .op(n19165) );
  nand2_1 U22749 ( .ip1(n19168), .ip2(n19165), .op(n18758) );
  buf_1 U22750 ( .ip(n24329), .op(n24180) );
  nand2_1 U22751 ( .ip1(\x[65][15] ), .ip2(n24180), .op(n18831) );
  nand2_1 U22752 ( .ip1(n18758), .ip2(n18831), .op(n18838) );
  inv_1 U22753 ( .ip(n18841), .op(n18759) );
  or2_1 U22754 ( .ip1(\x[66][12] ), .ip2(n18759), .op(n18761) );
  or2_1 U22755 ( .ip1(n24449), .ip2(n18759), .op(n18760) );
  nand2_1 U22756 ( .ip1(n18761), .ip2(n18760), .op(n19105) );
  nor2_1 U22757 ( .ip1(n24456), .ip2(\x[66][11] ), .op(n18790) );
  and2_1 U22758 ( .ip1(n24451), .ip2(\x[66][10] ), .op(n18788) );
  nand2_1 U22759 ( .ip1(\x[66][7] ), .ip2(n24461), .op(n18782) );
  nand2_1 U22760 ( .ip1(\x[66][8] ), .ip2(n24491), .op(n18781) );
  nand2_1 U22761 ( .ip1(\x[66][9] ), .ip2(n24269), .op(n18780) );
  and2_1 U22762 ( .ip1(n23283), .ip2(\x[66][5] ), .op(n18770) );
  inv_1 U22763 ( .ip(\x[66][3] ), .op(n18768) );
  inv_1 U22764 ( .ip(\x[66][1] ), .op(n18763) );
  nor2_1 U22765 ( .ip1(n22513), .ip2(n18763), .op(n18765) );
  inv_1 U22766 ( .ip(\x[66][0] ), .op(n18762) );
  not_ab_or_c_or_d U22767 ( .ip1(n24467), .ip2(n18763), .ip3(sig_in[0]), .ip4(
        n18762), .op(n18764) );
  not_ab_or_c_or_d U22768 ( .ip1(\x[66][2] ), .ip2(n24335), .ip3(n18765), 
        .ip4(n18764), .op(n18767) );
  nor2_1 U22769 ( .ip1(\x[66][2] ), .ip2(n24463), .op(n18766) );
  not_ab_or_c_or_d U22770 ( .ip1(n23251), .ip2(n18768), .ip3(n18767), .ip4(
        n18766), .op(n18769) );
  not_ab_or_c_or_d U22771 ( .ip1(\x[66][3] ), .ip2(n22795), .ip3(n18770), 
        .ip4(n18769), .op(n18774) );
  nand2_1 U22772 ( .ip1(\x[66][4] ), .ip2(n23721), .op(n18773) );
  not_ab_or_c_or_d U22773 ( .ip1(\x[66][5] ), .ip2(n23600), .ip3(\x[66][4] ), 
        .ip4(n24347), .op(n18772) );
  nor2_1 U22774 ( .ip1(\x[66][5] ), .ip2(n24119), .op(n18771) );
  not_ab_or_c_or_d U22775 ( .ip1(n18774), .ip2(n18773), .ip3(n18772), .ip4(
        n18771), .op(n18775) );
  nand2_1 U22776 ( .ip1(n18775), .ip2(\x[66][6] ), .op(n18778) );
  nor2_1 U22777 ( .ip1(\x[66][7] ), .ip2(n24142), .op(n18777) );
  nor2_1 U22778 ( .ip1(n18775), .ip2(\x[66][6] ), .op(n18776) );
  ab_or_c_or_d U22779 ( .ip1(sig_in[6]), .ip2(n18778), .ip3(n18777), .ip4(
        n18776), .op(n18779) );
  and4_1 U22780 ( .ip1(n18782), .ip2(n18781), .ip3(n18780), .ip4(n18779), .op(
        n18786) );
  nor2_1 U22781 ( .ip1(\x[66][10] ), .ip2(n20880), .op(n18785) );
  not_ab_or_c_or_d U22782 ( .ip1(\x[66][9] ), .ip2(n24043), .ip3(\x[66][8] ), 
        .ip4(n24358), .op(n18784) );
  nor2_1 U22783 ( .ip1(\x[66][9] ), .ip2(n24043), .op(n18783) );
  nor4_1 U22784 ( .ip1(n18786), .ip2(n18785), .ip3(n18784), .ip4(n18783), .op(
        n18787) );
  not_ab_or_c_or_d U22785 ( .ip1(\x[66][11] ), .ip2(n24371), .ip3(n18788), 
        .ip4(n18787), .op(n18789) );
  nor2_1 U22786 ( .ip1(n18790), .ip2(n18789), .op(n19113) );
  inv_1 U22787 ( .ip(n19113), .op(n18791) );
  nand2_1 U22788 ( .ip1(n19105), .ip2(n18791), .op(n18837) );
  nand2_1 U22789 ( .ip1(\x[65][10] ), .ip2(n23980), .op(n18818) );
  nor2_1 U22790 ( .ip1(\x[65][9] ), .ip2(n23981), .op(n18813) );
  inv_1 U22791 ( .ip(\x[65][8] ), .op(n18792) );
  nor3_1 U22792 ( .ip1(sig_in[8]), .ip2(n18813), .ip3(n18792), .op(n18816) );
  and2_1 U22793 ( .ip1(n24461), .ip2(\x[65][7] ), .op(n18810) );
  nor2_1 U22794 ( .ip1(n24347), .ip2(\x[65][4] ), .op(n18803) );
  inv_1 U22795 ( .ip(\x[65][3] ), .op(n18799) );
  nor2_1 U22796 ( .ip1(sig_in[3]), .ip2(n18799), .op(n18801) );
  inv_1 U22797 ( .ip(\x[65][1] ), .op(n18794) );
  nor2_1 U22798 ( .ip1(n22513), .ip2(n18794), .op(n18796) );
  inv_1 U22799 ( .ip(\x[65][0] ), .op(n18793) );
  not_ab_or_c_or_d U22800 ( .ip1(n24467), .ip2(n18794), .ip3(sig_in[0]), .ip4(
        n18793), .op(n18795) );
  not_ab_or_c_or_d U22801 ( .ip1(\x[65][2] ), .ip2(n24470), .ip3(n18796), 
        .ip4(n18795), .op(n18798) );
  nor2_1 U22802 ( .ip1(\x[65][2] ), .ip2(n24463), .op(n18797) );
  not_ab_or_c_or_d U22803 ( .ip1(n23251), .ip2(n18799), .ip3(n18798), .ip4(
        n18797), .op(n18800) );
  not_ab_or_c_or_d U22804 ( .ip1(\x[65][4] ), .ip2(n23860), .ip3(n18801), 
        .ip4(n18800), .op(n18802) );
  or2_1 U22805 ( .ip1(n18803), .ip2(n18802), .op(n18806) );
  nor2_1 U22806 ( .ip1(\x[65][6] ), .ip2(n23770), .op(n18805) );
  nor3_1 U22807 ( .ip1(n22833), .ip2(n18806), .ip3(n18805), .op(n18808) );
  inv_1 U22808 ( .ip(\x[65][5] ), .op(n18804) );
  not_ab_or_c_or_d U22809 ( .ip1(n18806), .ip2(n22833), .ip3(n18805), .ip4(
        n18804), .op(n18807) );
  or2_1 U22810 ( .ip1(n18808), .ip2(n18807), .op(n18809) );
  not_ab_or_c_or_d U22811 ( .ip1(\x[65][6] ), .ip2(n23770), .ip3(n18810), 
        .ip4(n18809), .op(n18814) );
  nor2_1 U22812 ( .ip1(\x[65][8] ), .ip2(n23971), .op(n18812) );
  nor2_1 U22813 ( .ip1(\x[65][7] ), .ip2(n24142), .op(n18811) );
  nor4_1 U22814 ( .ip1(n18814), .ip2(n18813), .ip3(n18812), .ip4(n18811), .op(
        n18815) );
  not_ab_or_c_or_d U22815 ( .ip1(\x[65][9] ), .ip2(n23981), .ip3(n18816), 
        .ip4(n18815), .op(n18817) );
  nand2_1 U22816 ( .ip1(n18818), .ip2(n18817), .op(n18824) );
  nor2_1 U22817 ( .ip1(\x[65][10] ), .ip2(n20880), .op(n18819) );
  or2_1 U22818 ( .ip1(sig_in[11]), .ip2(n18819), .op(n18822) );
  inv_1 U22819 ( .ip(\x[65][11] ), .op(n18820) );
  or2_1 U22820 ( .ip1(n18820), .ip2(n18819), .op(n18821) );
  nand2_1 U22821 ( .ip1(n18822), .ip2(n18821), .op(n18823) );
  nand2_1 U22822 ( .ip1(n18824), .ip2(n18823), .op(n18826) );
  nand2_1 U22823 ( .ip1(\x[65][11] ), .ip2(n24456), .op(n18825) );
  nand2_1 U22824 ( .ip1(n18826), .ip2(n18825), .op(n19163) );
  nor2_1 U22825 ( .ip1(\x[65][13] ), .ip2(n24235), .op(n18827) );
  or2_1 U22826 ( .ip1(n17845), .ip2(n18827), .op(n18830) );
  inv_1 U22827 ( .ip(\x[65][12] ), .op(n18828) );
  or2_1 U22828 ( .ip1(n18828), .ip2(n18827), .op(n18829) );
  nand2_1 U22829 ( .ip1(n18830), .ip2(n18829), .op(n19166) );
  inv_1 U22830 ( .ip(n18831), .op(n18832) );
  or2_1 U22831 ( .ip1(sig_in[14]), .ip2(n18832), .op(n18835) );
  inv_1 U22832 ( .ip(\x[65][14] ), .op(n18833) );
  or2_1 U22833 ( .ip1(n18833), .ip2(n18832), .op(n18834) );
  nand2_1 U22834 ( .ip1(n18835), .ip2(n18834), .op(n19172) );
  nand3_1 U22835 ( .ip1(n19163), .ip2(n19166), .ip3(n19172), .op(n18836) );
  nand3_1 U22836 ( .ip1(n18838), .ip2(n18837), .ip3(n18836), .op(n18839) );
  not_ab_or_c_or_d U22837 ( .ip1(n18841), .ip2(n18840), .ip3(n19104), .ip4(
        n18839), .op(n24657) );
  and2_1 U22838 ( .ip1(n23895), .ip2(\x[67][13] ), .op(n18842) );
  nor2_1 U22839 ( .ip1(\x[67][15] ), .ip2(n23143), .op(n19108) );
  not_ab_or_c_or_d U22840 ( .ip1(\x[67][14] ), .ip2(n24185), .ip3(n18842), 
        .ip4(n19108), .op(n19112) );
  nand2_1 U22841 ( .ip1(\x[67][12] ), .ip2(n24233), .op(n18843) );
  nand2_1 U22842 ( .ip1(n19112), .ip2(n18843), .op(n19101) );
  nand2_1 U22843 ( .ip1(\x[67][15] ), .ip2(n24180), .op(n18932) );
  nor2_1 U22844 ( .ip1(\x[68][14] ), .ip2(n24230), .op(n18888) );
  inv_1 U22845 ( .ip(\x[68][12] ), .op(n18882) );
  inv_1 U22846 ( .ip(\x[68][9] ), .op(n18865) );
  nand2_1 U22847 ( .ip1(n21171), .ip2(n18865), .op(n18871) );
  inv_1 U22848 ( .ip(\x[68][10] ), .op(n18872) );
  not_ab_or_c_or_d U22849 ( .ip1(\x[68][9] ), .ip2(n23981), .ip3(\x[68][8] ), 
        .ip4(n24358), .op(n18869) );
  inv_1 U22850 ( .ip(\x[68][7] ), .op(n18862) );
  nor2_1 U22851 ( .ip1(n17732), .ip2(n18862), .op(n18860) );
  inv_1 U22852 ( .ip(\x[68][3] ), .op(n18850) );
  inv_1 U22853 ( .ip(\x[68][1] ), .op(n18845) );
  nor2_1 U22854 ( .ip1(n22513), .ip2(n18845), .op(n18847) );
  inv_1 U22855 ( .ip(\x[68][0] ), .op(n18844) );
  not_ab_or_c_or_d U22856 ( .ip1(n24467), .ip2(n18845), .ip3(sig_in[0]), .ip4(
        n18844), .op(n18846) );
  not_ab_or_c_or_d U22857 ( .ip1(\x[68][2] ), .ip2(n24335), .ip3(n18847), 
        .ip4(n18846), .op(n18849) );
  buf_1 U22858 ( .ip(n24107), .op(n23717) );
  nor2_1 U22859 ( .ip1(\x[68][2] ), .ip2(n23717), .op(n18848) );
  not_ab_or_c_or_d U22860 ( .ip1(n24251), .ip2(n18850), .ip3(n18849), .ip4(
        n18848), .op(n18854) );
  nand2_1 U22861 ( .ip1(\x[68][5] ), .ip2(n24350), .op(n18852) );
  nand2_1 U22862 ( .ip1(\x[68][4] ), .ip2(n23721), .op(n18851) );
  nand2_1 U22863 ( .ip1(n18852), .ip2(n18851), .op(n18853) );
  not_ab_or_c_or_d U22864 ( .ip1(\x[68][3] ), .ip2(n22795), .ip3(n18854), 
        .ip4(n18853), .op(n18858) );
  nor2_1 U22865 ( .ip1(\x[68][6] ), .ip2(n23770), .op(n18857) );
  nor2_1 U22866 ( .ip1(\x[68][5] ), .ip2(n24350), .op(n18856) );
  not_ab_or_c_or_d U22867 ( .ip1(\x[68][5] ), .ip2(n23600), .ip3(\x[68][4] ), 
        .ip4(n24347), .op(n18855) );
  nor4_1 U22868 ( .ip1(n18858), .ip2(n18857), .ip3(n18856), .ip4(n18855), .op(
        n18859) );
  not_ab_or_c_or_d U22869 ( .ip1(\x[68][6] ), .ip2(n24355), .ip3(n18860), 
        .ip4(n18859), .op(n18861) );
  or2_1 U22870 ( .ip1(sig_in[7]), .ip2(n18861), .op(n18864) );
  or2_1 U22871 ( .ip1(n18862), .ip2(n18861), .op(n18863) );
  nand2_1 U22872 ( .ip1(n18864), .ip2(n18863), .op(n18867) );
  nor2_1 U22873 ( .ip1(n21171), .ip2(n18865), .op(n18866) );
  not_ab_or_c_or_d U22874 ( .ip1(\x[68][8] ), .ip2(n24491), .ip3(n18867), 
        .ip4(n18866), .op(n18868) );
  not_ab_or_c_or_d U22875 ( .ip1(sig_in[10]), .ip2(n18872), .ip3(n18869), 
        .ip4(n18868), .op(n18870) );
  nand2_1 U22876 ( .ip1(n18871), .ip2(n18870), .op(n18877) );
  nor2_1 U22877 ( .ip1(sig_in[10]), .ip2(n18872), .op(n18873) );
  or2_1 U22878 ( .ip1(\x[68][11] ), .ip2(n18873), .op(n18875) );
  or2_1 U22879 ( .ip1(n24456), .ip2(n18873), .op(n18874) );
  nand2_1 U22880 ( .ip1(n18875), .ip2(n18874), .op(n18876) );
  nand2_1 U22881 ( .ip1(n18877), .ip2(n18876), .op(n18879) );
  or2_1 U22882 ( .ip1(n24136), .ip2(\x[68][11] ), .op(n18878) );
  nand2_1 U22883 ( .ip1(n18879), .ip2(n18878), .op(n18881) );
  nor2_1 U22884 ( .ip1(\x[68][13] ), .ip2(n24137), .op(n18880) );
  not_ab_or_c_or_d U22885 ( .ip1(n17845), .ip2(n18882), .ip3(n18881), .ip4(
        n18880), .op(n18886) );
  nand2_1 U22886 ( .ip1(\x[68][13] ), .ip2(n24081), .op(n18884) );
  nand2_1 U22887 ( .ip1(\x[68][12] ), .ip2(n24233), .op(n18883) );
  nand2_1 U22888 ( .ip1(n18884), .ip2(n18883), .op(n18885) );
  not_ab_or_c_or_d U22889 ( .ip1(\x[68][14] ), .ip2(n24230), .ip3(n18886), 
        .ip4(n18885), .op(n18887) );
  not_ab_or_c_or_d U22890 ( .ip1(\x[68][15] ), .ip2(n24384), .ip3(n18888), 
        .ip4(n18887), .op(n18890) );
  nor2_1 U22891 ( .ip1(\x[68][15] ), .ip2(n23143), .op(n18889) );
  nor2_1 U22892 ( .ip1(n18890), .ip2(n18889), .op(n19096) );
  inv_1 U22893 ( .ip(\x[67][11] ), .op(n18924) );
  and2_1 U22894 ( .ip1(n24451), .ip2(\x[67][10] ), .op(n18921) );
  inv_1 U22895 ( .ip(\x[67][7] ), .op(n18914) );
  inv_1 U22896 ( .ip(\x[67][6] ), .op(n18906) );
  nor2_1 U22897 ( .ip1(sig_in[6]), .ip2(n18906), .op(n18904) );
  inv_1 U22898 ( .ip(\x[67][4] ), .op(n18902) );
  nor2_1 U22899 ( .ip1(n24462), .ip2(n18902), .op(n18899) );
  inv_1 U22900 ( .ip(\x[67][3] ), .op(n18897) );
  inv_1 U22901 ( .ip(\x[67][1] ), .op(n18892) );
  nor2_1 U22902 ( .ip1(n24467), .ip2(n18892), .op(n18894) );
  inv_1 U22903 ( .ip(\x[67][0] ), .op(n18891) );
  not_ab_or_c_or_d U22904 ( .ip1(sig_in[1]), .ip2(n18892), .ip3(sig_in[0]), 
        .ip4(n18891), .op(n18893) );
  not_ab_or_c_or_d U22905 ( .ip1(\x[67][2] ), .ip2(n23659), .ip3(n18894), 
        .ip4(n18893), .op(n18896) );
  nor2_1 U22906 ( .ip1(\x[67][2] ), .ip2(n24463), .op(n18895) );
  not_ab_or_c_or_d U22907 ( .ip1(n23251), .ip2(n18897), .ip3(n18896), .ip4(
        n18895), .op(n18898) );
  not_ab_or_c_or_d U22908 ( .ip1(\x[67][3] ), .ip2(n22795), .ip3(n18899), 
        .ip4(n18898), .op(n18901) );
  nor2_1 U22909 ( .ip1(\x[67][5] ), .ip2(n23283), .op(n18900) );
  not_ab_or_c_or_d U22910 ( .ip1(sig_in[4]), .ip2(n18902), .ip3(n18901), .ip4(
        n18900), .op(n18903) );
  not_ab_or_c_or_d U22911 ( .ip1(\x[67][5] ), .ip2(n23600), .ip3(n18904), 
        .ip4(n18903), .op(n18905) );
  or2_1 U22912 ( .ip1(sig_in[6]), .ip2(n18905), .op(n18908) );
  or2_1 U22913 ( .ip1(n18906), .ip2(n18905), .op(n18907) );
  nand2_1 U22914 ( .ip1(n18908), .ip2(n18907), .op(n18909) );
  or2_1 U22915 ( .ip1(\x[67][7] ), .ip2(n18909), .op(n18911) );
  or2_1 U22916 ( .ip1(n24142), .ip2(n18909), .op(n18910) );
  nand2_1 U22917 ( .ip1(n18911), .ip2(n18910), .op(n18913) );
  nor2_1 U22918 ( .ip1(\x[67][8] ), .ip2(n23971), .op(n18912) );
  not_ab_or_c_or_d U22919 ( .ip1(sig_in[7]), .ip2(n18914), .ip3(n18913), .ip4(
        n18912), .op(n18915) );
  or2_1 U22920 ( .ip1(\x[67][8] ), .ip2(n18915), .op(n18917) );
  or2_1 U22921 ( .ip1(n24491), .ip2(n18915), .op(n18916) );
  nand2_1 U22922 ( .ip1(n18917), .ip2(n18916), .op(n18919) );
  nor2_1 U22923 ( .ip1(\x[67][9] ), .ip2(n24269), .op(n18918) );
  nor2_1 U22924 ( .ip1(n18919), .ip2(n18918), .op(n18920) );
  not_ab_or_c_or_d U22925 ( .ip1(\x[67][9] ), .ip2(n23981), .ip3(n18921), 
        .ip4(n18920), .op(n18923) );
  nor2_1 U22926 ( .ip1(\x[67][10] ), .ip2(n20880), .op(n18922) );
  not_ab_or_c_or_d U22927 ( .ip1(sig_in[11]), .ip2(n18924), .ip3(n18923), 
        .ip4(n18922), .op(n18925) );
  or2_1 U22928 ( .ip1(\x[67][11] ), .ip2(n18925), .op(n18927) );
  or2_1 U22929 ( .ip1(n24136), .ip2(n18925), .op(n18926) );
  nand2_1 U22930 ( .ip1(n18927), .ip2(n18926), .op(n19103) );
  nor2_1 U22931 ( .ip1(\x[67][13] ), .ip2(n24376), .op(n18929) );
  nor2_1 U22932 ( .ip1(\x[67][12] ), .ip2(n24449), .op(n18928) );
  or2_1 U22933 ( .ip1(n18929), .ip2(n18928), .op(n19111) );
  or2_1 U22934 ( .ip1(n24185), .ip2(\x[67][14] ), .op(n18930) );
  nand2_1 U22935 ( .ip1(n18932), .ip2(n18930), .op(n19106) );
  nor3_1 U22936 ( .ip1(n19103), .ip2(n19111), .ip3(n19106), .op(n18931) );
  not_ab_or_c_or_d U22937 ( .ip1(n19101), .ip2(n18932), .ip3(n19096), .ip4(
        n18931), .op(n24660) );
  nand2_1 U22938 ( .ip1(\x[70][15] ), .ip2(n24186), .op(n19018) );
  and2_1 U22939 ( .ip1(n23895), .ip2(\x[70][13] ), .op(n18933) );
  nor2_1 U22940 ( .ip1(\x[70][15] ), .ip2(n23143), .op(n19019) );
  not_ab_or_c_or_d U22941 ( .ip1(\x[70][14] ), .ip2(n24185), .ip3(n18933), 
        .ip4(n19019), .op(n19038) );
  nand2_1 U22942 ( .ip1(\x[70][12] ), .ip2(n24449), .op(n18934) );
  nand2_1 U22943 ( .ip1(n19038), .ip2(n18934), .op(n19033) );
  and2_1 U22944 ( .ip1(n24451), .ip2(\x[70][10] ), .op(n18935) );
  and2_1 U22945 ( .ip1(n24371), .ip2(\x[70][11] ), .op(n18939) );
  not_ab_or_c_or_d U22946 ( .ip1(\x[70][9] ), .ip2(n23981), .ip3(n18935), 
        .ip4(n18939), .op(n19024) );
  inv_1 U22947 ( .ip(\x[70][8] ), .op(n18943) );
  nor2_1 U22948 ( .ip1(n24455), .ip2(\x[70][9] ), .op(n18942) );
  or3_1 U22949 ( .ip1(n23779), .ip2(n18943), .ip3(n18942), .op(n18936) );
  nand2_1 U22950 ( .ip1(n19024), .ip2(n18936), .op(n18941) );
  nor2_1 U22951 ( .ip1(\x[70][11] ), .ip2(n24456), .op(n18938) );
  nor2_1 U22952 ( .ip1(\x[70][10] ), .ip2(n20880), .op(n18937) );
  nor2_1 U22953 ( .ip1(n18938), .ip2(n18937), .op(n18966) );
  nor2_1 U22954 ( .ip1(n18939), .ip2(n18966), .op(n19030) );
  inv_1 U22955 ( .ip(n19030), .op(n18940) );
  nand2_1 U22956 ( .ip1(n18941), .ip2(n18940), .op(n18971) );
  or2_1 U22957 ( .ip1(n23779), .ip2(n18942), .op(n18945) );
  or2_1 U22958 ( .ip1(n18943), .ip2(n18942), .op(n18944) );
  nand2_1 U22959 ( .ip1(n18945), .ip2(n18944), .op(n19028) );
  inv_1 U22960 ( .ip(\x[70][7] ), .op(n18962) );
  nor2_1 U22961 ( .ip1(n18962), .ip2(n17732), .op(n18964) );
  and2_1 U22962 ( .ip1(n24485), .ip2(\x[70][6] ), .op(n18959) );
  inv_1 U22963 ( .ip(\x[70][4] ), .op(n18957) );
  nor2_1 U22964 ( .ip1(n24462), .ip2(n18957), .op(n18954) );
  inv_1 U22965 ( .ip(\x[70][3] ), .op(n18952) );
  inv_1 U22966 ( .ip(\x[70][1] ), .op(n18947) );
  nor2_1 U22967 ( .ip1(n22513), .ip2(n18947), .op(n18949) );
  inv_1 U22968 ( .ip(\x[70][0] ), .op(n18946) );
  not_ab_or_c_or_d U22969 ( .ip1(sig_in[1]), .ip2(n18947), .ip3(n23195), .ip4(
        n18946), .op(n18948) );
  not_ab_or_c_or_d U22970 ( .ip1(\x[70][2] ), .ip2(n24470), .ip3(n18949), 
        .ip4(n18948), .op(n18951) );
  nor2_1 U22971 ( .ip1(\x[70][2] ), .ip2(n24463), .op(n18950) );
  not_ab_or_c_or_d U22972 ( .ip1(n24251), .ip2(n18952), .ip3(n18951), .ip4(
        n18950), .op(n18953) );
  not_ab_or_c_or_d U22973 ( .ip1(\x[70][3] ), .ip2(n22795), .ip3(n18954), 
        .ip4(n18953), .op(n18956) );
  nor2_1 U22974 ( .ip1(\x[70][5] ), .ip2(n24119), .op(n18955) );
  not_ab_or_c_or_d U22975 ( .ip1(sig_in[4]), .ip2(n18957), .ip3(n18956), .ip4(
        n18955), .op(n18958) );
  not_ab_or_c_or_d U22976 ( .ip1(\x[70][5] ), .ip2(n23600), .ip3(n18959), 
        .ip4(n18958), .op(n18961) );
  nor2_1 U22977 ( .ip1(\x[70][6] ), .ip2(n24485), .op(n18960) );
  not_ab_or_c_or_d U22978 ( .ip1(sig_in[7]), .ip2(n18962), .ip3(n18961), .ip4(
        n18960), .op(n18963) );
  nor2_1 U22979 ( .ip1(n18964), .ip2(n18963), .op(n19031) );
  inv_1 U22980 ( .ip(n19031), .op(n18965) );
  nand3_1 U22981 ( .ip1(n18966), .ip2(n19028), .ip3(n18965), .op(n18970) );
  or2_1 U22982 ( .ip1(n24382), .ip2(\x[70][14] ), .op(n18967) );
  nand2_1 U22983 ( .ip1(n19018), .ip2(n18967), .op(n19086) );
  nor2_1 U22984 ( .ip1(\x[70][13] ), .ip2(n24081), .op(n18969) );
  nor2_1 U22985 ( .ip1(\x[70][12] ), .ip2(n24079), .op(n18968) );
  or2_1 U22986 ( .ip1(n18969), .ip2(n18968), .op(n19037) );
  not_ab_or_c_or_d U22987 ( .ip1(n18971), .ip2(n18970), .ip3(n19086), .ip4(
        n19037), .op(n19017) );
  inv_1 U22988 ( .ip(\x[71][9] ), .op(n18972) );
  nand2_1 U22989 ( .ip1(n21171), .ip2(n18972), .op(n18997) );
  nor2_1 U22990 ( .ip1(n21171), .ip2(n18972), .op(n18991) );
  inv_1 U22991 ( .ip(\x[71][6] ), .op(n18989) );
  nor2_1 U22992 ( .ip1(sig_in[6]), .ip2(n18989), .op(n18986) );
  inv_1 U22993 ( .ip(\x[71][4] ), .op(n18984) );
  nor2_1 U22994 ( .ip1(n24462), .ip2(n18984), .op(n18981) );
  inv_1 U22995 ( .ip(\x[71][3] ), .op(n18979) );
  nor2_1 U22996 ( .ip1(\x[71][2] ), .ip2(n24463), .op(n18978) );
  inv_1 U22997 ( .ip(\x[71][1] ), .op(n18974) );
  nor2_1 U22998 ( .ip1(n22513), .ip2(n18974), .op(n18976) );
  inv_1 U22999 ( .ip(\x[71][0] ), .op(n18973) );
  not_ab_or_c_or_d U23000 ( .ip1(sig_in[1]), .ip2(n18974), .ip3(sig_in[0]), 
        .ip4(n18973), .op(n18975) );
  not_ab_or_c_or_d U23001 ( .ip1(\x[71][2] ), .ip2(n24335), .ip3(n18976), 
        .ip4(n18975), .op(n18977) );
  not_ab_or_c_or_d U23002 ( .ip1(n24251), .ip2(n18979), .ip3(n18978), .ip4(
        n18977), .op(n18980) );
  not_ab_or_c_or_d U23003 ( .ip1(\x[71][3] ), .ip2(n22795), .ip3(n18981), 
        .ip4(n18980), .op(n18983) );
  nor2_1 U23004 ( .ip1(\x[71][5] ), .ip2(n24350), .op(n18982) );
  not_ab_or_c_or_d U23005 ( .ip1(sig_in[4]), .ip2(n18984), .ip3(n18983), .ip4(
        n18982), .op(n18985) );
  not_ab_or_c_or_d U23006 ( .ip1(\x[71][5] ), .ip2(n23600), .ip3(n18986), 
        .ip4(n18985), .op(n18988) );
  nor2_1 U23007 ( .ip1(\x[71][7] ), .ip2(n24142), .op(n18987) );
  not_ab_or_c_or_d U23008 ( .ip1(sig_in[6]), .ip2(n18989), .ip3(n18988), .ip4(
        n18987), .op(n18990) );
  not_ab_or_c_or_d U23009 ( .ip1(\x[71][7] ), .ip2(n24142), .ip3(n18991), 
        .ip4(n18990), .op(n18995) );
  nand2_1 U23010 ( .ip1(\x[71][8] ), .ip2(n23971), .op(n18994) );
  nor2_1 U23011 ( .ip1(\x[71][10] ), .ip2(n20880), .op(n18993) );
  not_ab_or_c_or_d U23012 ( .ip1(\x[71][9] ), .ip2(n23981), .ip3(\x[71][8] ), 
        .ip4(n24358), .op(n18992) );
  not_ab_or_c_or_d U23013 ( .ip1(n18995), .ip2(n18994), .ip3(n18993), .ip4(
        n18992), .op(n18996) );
  nand2_1 U23014 ( .ip1(n18997), .ip2(n18996), .op(n19002) );
  buf_1 U23015 ( .ip(n24370), .op(n23146) );
  and2_1 U23016 ( .ip1(n23146), .ip2(\x[71][10] ), .op(n18998) );
  or2_1 U23017 ( .ip1(\x[71][11] ), .ip2(n18998), .op(n19000) );
  or2_1 U23018 ( .ip1(n24136), .ip2(n18998), .op(n18999) );
  nand2_1 U23019 ( .ip1(n19000), .ip2(n18999), .op(n19001) );
  nand2_1 U23020 ( .ip1(n19002), .ip2(n19001), .op(n19004) );
  or2_1 U23021 ( .ip1(n21793), .ip2(\x[71][11] ), .op(n19003) );
  and2_1 U23022 ( .ip1(n19004), .ip2(n19003), .op(n20055) );
  inv_1 U23023 ( .ip(\x[71][12] ), .op(n19006) );
  nor2_1 U23024 ( .ip1(n19006), .ip2(n17845), .op(n20053) );
  or2_1 U23025 ( .ip1(n20055), .ip2(n20053), .op(n19009) );
  nor2_1 U23026 ( .ip1(\x[71][13] ), .ip2(n23895), .op(n19005) );
  or2_1 U23027 ( .ip1(n17845), .ip2(n19005), .op(n19008) );
  or2_1 U23028 ( .ip1(n19006), .ip2(n19005), .op(n19007) );
  nand2_1 U23029 ( .ip1(n19008), .ip2(n19007), .op(n20056) );
  nand2_1 U23030 ( .ip1(n19009), .ip2(n20056), .op(n19011) );
  and2_1 U23031 ( .ip1(n24332), .ip2(\x[71][13] ), .op(n20054) );
  nor2_1 U23032 ( .ip1(\x[71][15] ), .ip2(n23143), .op(n20059) );
  not_ab_or_c_or_d U23033 ( .ip1(\x[71][14] ), .ip2(n24185), .ip3(n20054), 
        .ip4(n20059), .op(n19010) );
  nand2_1 U23034 ( .ip1(n19011), .ip2(n19010), .op(n19015) );
  inv_1 U23035 ( .ip(n20059), .op(n19013) );
  nand2_1 U23036 ( .ip1(\x[71][15] ), .ip2(n24180), .op(n20062) );
  or2_1 U23037 ( .ip1(n24185), .ip2(\x[71][14] ), .op(n19012) );
  nand2_1 U23038 ( .ip1(n20062), .ip2(n19012), .op(n20057) );
  nand2_1 U23039 ( .ip1(n19013), .ip2(n20057), .op(n19014) );
  nand2_1 U23040 ( .ip1(n19015), .ip2(n19014), .op(n19016) );
  not_ab_or_c_or_d U23041 ( .ip1(n19018), .ip2(n19033), .ip3(n19017), .ip4(
        n19016), .op(n27536) );
  inv_1 U23042 ( .ip(n19019), .op(n19085) );
  nor2_1 U23043 ( .ip1(\x[69][15] ), .ip2(n23143), .op(n19093) );
  inv_1 U23044 ( .ip(\x[69][14] ), .op(n19044) );
  nor2_1 U23045 ( .ip1(sig_in[14]), .ip2(n19044), .op(n19021) );
  and2_1 U23046 ( .ip1(n24332), .ip2(\x[69][13] ), .op(n19020) );
  nor2_1 U23047 ( .ip1(n19021), .ip2(n19020), .op(n19091) );
  and2_1 U23048 ( .ip1(n24186), .ip2(\x[69][15] ), .op(n19043) );
  or2_1 U23049 ( .ip1(n19091), .ip2(n19043), .op(n19023) );
  nand2_1 U23050 ( .ip1(\x[69][12] ), .ip2(n24233), .op(n19089) );
  or2_1 U23051 ( .ip1(n19089), .ip2(n19043), .op(n19022) );
  nand2_1 U23052 ( .ip1(n19023), .ip2(n19022), .op(n19036) );
  inv_1 U23053 ( .ip(n19024), .op(n19027) );
  or2_1 U23054 ( .ip1(\x[70][8] ), .ip2(n19027), .op(n19026) );
  or2_1 U23055 ( .ip1(n24491), .ip2(n19027), .op(n19025) );
  nand2_1 U23056 ( .ip1(n19026), .ip2(n19025), .op(n19032) );
  nor2_1 U23057 ( .ip1(n19028), .ip2(n19027), .op(n19029) );
  not_ab_or_c_or_d U23058 ( .ip1(n19032), .ip2(n19031), .ip3(n19030), .ip4(
        n19029), .op(n19034) );
  nor2_1 U23059 ( .ip1(n19034), .ip2(n19033), .op(n19035) );
  not_ab_or_c_or_d U23060 ( .ip1(n19038), .ip2(n19037), .ip3(n19036), .ip4(
        n19035), .op(n19083) );
  nor2_1 U23061 ( .ip1(\x[69][13] ), .ip2(n24137), .op(n19039) );
  or2_1 U23062 ( .ip1(sig_in[12]), .ip2(n19039), .op(n19042) );
  inv_1 U23063 ( .ip(\x[69][12] ), .op(n19040) );
  or2_1 U23064 ( .ip1(n19040), .ip2(n19039), .op(n19041) );
  nand2_1 U23065 ( .ip1(n19042), .ip2(n19041), .op(n19095) );
  or2_1 U23066 ( .ip1(sig_in[14]), .ip2(n19043), .op(n19046) );
  or2_1 U23067 ( .ip1(n19044), .ip2(n19043), .op(n19045) );
  nand2_1 U23068 ( .ip1(n19046), .ip2(n19045), .op(n19087) );
  nor2_1 U23069 ( .ip1(\x[69][10] ), .ip2(n20880), .op(n19047) );
  or2_1 U23070 ( .ip1(sig_in[11]), .ip2(n19047), .op(n19050) );
  inv_1 U23071 ( .ip(\x[69][11] ), .op(n19048) );
  or2_1 U23072 ( .ip1(n19048), .ip2(n19047), .op(n19049) );
  nand2_1 U23073 ( .ip1(n19050), .ip2(n19049), .op(n19079) );
  inv_1 U23074 ( .ip(\x[69][7] ), .op(n19068) );
  nor2_1 U23075 ( .ip1(n19068), .ip2(n17732), .op(n19070) );
  nor2_1 U23076 ( .ip1(\x[69][6] ), .ip2(n23770), .op(n19067) );
  inv_1 U23077 ( .ip(n23251), .op(n22525) );
  and2_1 U23078 ( .ip1(n24107), .ip2(\x[69][2] ), .op(n19056) );
  nand2_1 U23079 ( .ip1(\x[69][1] ), .ip2(n21685), .op(n19054) );
  nand2_1 U23080 ( .ip1(\x[69][0] ), .ip2(n24143), .op(n19053) );
  nor2_1 U23081 ( .ip1(\x[69][2] ), .ip2(n24463), .op(n19052) );
  nor2_1 U23082 ( .ip1(\x[69][1] ), .ip2(n21685), .op(n19051) );
  not_ab_or_c_or_d U23083 ( .ip1(n19054), .ip2(n19053), .ip3(n19052), .ip4(
        n19051), .op(n19055) );
  not_ab_or_c_or_d U23084 ( .ip1(\x[69][3] ), .ip2(n22525), .ip3(n19056), 
        .ip4(n19055), .op(n19059) );
  nor2_1 U23085 ( .ip1(\x[69][5] ), .ip2(n24482), .op(n19060) );
  nor2_1 U23086 ( .ip1(\x[69][4] ), .ip2(n24347), .op(n19058) );
  nor2_1 U23087 ( .ip1(\x[69][3] ), .ip2(n24342), .op(n19057) );
  nor4_1 U23088 ( .ip1(n19059), .ip2(n19060), .ip3(n19058), .ip4(n19057), .op(
        n19065) );
  inv_1 U23089 ( .ip(n19060), .op(n19061) );
  nand3_1 U23090 ( .ip1(n23721), .ip2(\x[69][4] ), .ip3(n19061), .op(n19063)
         );
  nand2_1 U23091 ( .ip1(\x[69][6] ), .ip2(n24485), .op(n19062) );
  nand2_1 U23092 ( .ip1(n19063), .ip2(n19062), .op(n19064) );
  not_ab_or_c_or_d U23093 ( .ip1(\x[69][5] ), .ip2(n23600), .ip3(n19065), 
        .ip4(n19064), .op(n19066) );
  not_ab_or_c_or_d U23094 ( .ip1(sig_in[7]), .ip2(n19068), .ip3(n19067), .ip4(
        n19066), .op(n19069) );
  or2_1 U23095 ( .ip1(n19070), .ip2(n19069), .op(n19071) );
  nand2_1 U23096 ( .ip1(n19071), .ip2(\x[69][8] ), .op(n19074) );
  nor2_1 U23097 ( .ip1(\x[69][9] ), .ip2(n24164), .op(n19073) );
  nor2_1 U23098 ( .ip1(n19071), .ip2(\x[69][8] ), .op(n19072) );
  ab_or_c_or_d U23099 ( .ip1(n23779), .ip2(n19074), .ip3(n19073), .ip4(n19072), 
        .op(n19077) );
  nand2_1 U23100 ( .ip1(\x[69][10] ), .ip2(n23980), .op(n19076) );
  nand2_1 U23101 ( .ip1(\x[69][9] ), .ip2(n24164), .op(n19075) );
  nand3_1 U23102 ( .ip1(n19077), .ip2(n19076), .ip3(n19075), .op(n19078) );
  nand2_1 U23103 ( .ip1(n19079), .ip2(n19078), .op(n19081) );
  nand2_1 U23104 ( .ip1(\x[69][11] ), .ip2(n24456), .op(n19080) );
  nand2_1 U23105 ( .ip1(n19081), .ip2(n19080), .op(n19088) );
  nand3_1 U23106 ( .ip1(n19095), .ip2(n19087), .ip3(n19088), .op(n19082) );
  nand2_1 U23107 ( .ip1(n19083), .ip2(n19082), .op(n19084) );
  not_ab_or_c_or_d U23108 ( .ip1(n19086), .ip2(n19085), .ip3(n19093), .ip4(
        n19084), .op(n27535) );
  nor2_1 U23109 ( .ip1(n27536), .ip2(n27535), .op(n24663) );
  inv_1 U23110 ( .ip(n19093), .op(n19100) );
  inv_1 U23111 ( .ip(n19087), .op(n19099) );
  inv_1 U23112 ( .ip(n19088), .op(n19090) );
  nand2_1 U23113 ( .ip1(n19090), .ip2(n19089), .op(n19094) );
  inv_1 U23114 ( .ip(n19091), .op(n19092) );
  not_ab_or_c_or_d U23115 ( .ip1(n19095), .ip2(n19094), .ip3(n19093), .ip4(
        n19092), .op(n19098) );
  inv_1 U23116 ( .ip(n19096), .op(n19097) );
  ab_or_c_or_d U23117 ( .ip1(n19100), .ip2(n19099), .ip3(n19098), .ip4(n19097), 
        .op(n24665) );
  nand2_1 U23118 ( .ip1(n24663), .ip2(n24665), .op(n24661) );
  nor2_1 U23119 ( .ip1(n24660), .ip2(n24661), .op(n24654) );
  inv_1 U23120 ( .ip(n19101), .op(n19102) );
  nand2_1 U23121 ( .ip1(n19103), .ip2(n19102), .op(n19118) );
  nor2_1 U23122 ( .ip1(n19105), .ip2(n19104), .op(n19110) );
  inv_1 U23123 ( .ip(n19106), .op(n19107) );
  nor2_1 U23124 ( .ip1(n19108), .ip2(n19107), .op(n19109) );
  not_ab_or_c_or_d U23125 ( .ip1(n19112), .ip2(n19111), .ip3(n19110), .ip4(
        n19109), .op(n19117) );
  nand3_1 U23126 ( .ip1(n19115), .ip2(n19114), .ip3(n19113), .op(n19116) );
  nand3_1 U23127 ( .ip1(n19118), .ip2(n19117), .ip3(n19116), .op(n24656) );
  nand2_1 U23128 ( .ip1(n24654), .ip2(n24656), .op(n24658) );
  nor2_1 U23129 ( .ip1(n24657), .ip2(n24658), .op(n24672) );
  inv_1 U23130 ( .ip(\x[64][12] ), .op(n19170) );
  nor2_1 U23131 ( .ip1(\x[64][13] ), .ip2(n24376), .op(n19121) );
  or2_1 U23132 ( .ip1(n24382), .ip2(\x[64][14] ), .op(n19120) );
  nand2_1 U23133 ( .ip1(\x[64][15] ), .ip2(n24180), .op(n19119) );
  nand2_1 U23134 ( .ip1(n19120), .ip2(n19119), .op(n19171) );
  not_ab_or_c_or_d U23135 ( .ip1(sig_in[12]), .ip2(n19170), .ip3(n19121), 
        .ip4(n19171), .op(n19258) );
  nor2_1 U23136 ( .ip1(\x[64][15] ), .ip2(n23143), .op(n19159) );
  or2_1 U23137 ( .ip1(n19258), .ip2(n19159), .op(n19162) );
  inv_1 U23138 ( .ip(\x[64][9] ), .op(n19123) );
  nor2_1 U23139 ( .ip1(\x[64][10] ), .ip2(n20880), .op(n19122) );
  nor2_1 U23140 ( .ip1(\x[64][11] ), .ip2(n24371), .op(n19152) );
  not_ab_or_c_or_d U23141 ( .ip1(n21171), .ip2(n19123), .ip3(n19122), .ip4(
        n19152), .op(n19149) );
  inv_1 U23142 ( .ip(\x[64][7] ), .op(n19144) );
  nor2_1 U23143 ( .ip1(n17732), .ip2(n19144), .op(n19141) );
  nor2_1 U23144 ( .ip1(n24347), .ip2(\x[64][4] ), .op(n19134) );
  inv_1 U23145 ( .ip(\x[64][3] ), .op(n19130) );
  nor2_1 U23146 ( .ip1(sig_in[3]), .ip2(n19130), .op(n19132) );
  inv_1 U23147 ( .ip(\x[64][1] ), .op(n19125) );
  nor2_1 U23148 ( .ip1(n22513), .ip2(n19125), .op(n19127) );
  inv_1 U23149 ( .ip(\x[64][0] ), .op(n19124) );
  not_ab_or_c_or_d U23150 ( .ip1(n24464), .ip2(n19125), .ip3(n23195), .ip4(
        n19124), .op(n19126) );
  not_ab_or_c_or_d U23151 ( .ip1(\x[64][2] ), .ip2(n23659), .ip3(n19127), 
        .ip4(n19126), .op(n19129) );
  nor2_1 U23152 ( .ip1(\x[64][2] ), .ip2(n24463), .op(n19128) );
  not_ab_or_c_or_d U23153 ( .ip1(n23251), .ip2(n19130), .ip3(n19129), .ip4(
        n19128), .op(n19131) );
  not_ab_or_c_or_d U23154 ( .ip1(\x[64][4] ), .ip2(n23860), .ip3(n19132), 
        .ip4(n19131), .op(n19133) );
  or2_1 U23155 ( .ip1(n19134), .ip2(n19133), .op(n19137) );
  nor2_1 U23156 ( .ip1(\x[64][6] ), .ip2(n23509), .op(n19136) );
  nor3_1 U23157 ( .ip1(n22833), .ip2(n19137), .ip3(n19136), .op(n19139) );
  inv_1 U23158 ( .ip(\x[64][5] ), .op(n19135) );
  not_ab_or_c_or_d U23159 ( .ip1(n19137), .ip2(n22833), .ip3(n19136), .ip4(
        n19135), .op(n19138) );
  or2_1 U23160 ( .ip1(n19139), .ip2(n19138), .op(n19140) );
  not_ab_or_c_or_d U23161 ( .ip1(\x[64][6] ), .ip2(n23509), .ip3(n19141), 
        .ip4(n19140), .op(n19143) );
  nor2_1 U23162 ( .ip1(\x[64][8] ), .ip2(n23971), .op(n19142) );
  ab_or_c_or_d U23163 ( .ip1(sig_in[7]), .ip2(n19144), .ip3(n19143), .ip4(
        n19142), .op(n19147) );
  nand2_1 U23164 ( .ip1(\x[64][8] ), .ip2(n23804), .op(n19146) );
  nand2_1 U23165 ( .ip1(\x[64][9] ), .ip2(n24164), .op(n19145) );
  nand3_1 U23166 ( .ip1(n19147), .ip2(n19146), .ip3(n19145), .op(n19148) );
  nand2_1 U23167 ( .ip1(n19149), .ip2(n19148), .op(n19158) );
  nand2_1 U23168 ( .ip1(n21793), .ip2(\x[64][11] ), .op(n19151) );
  nand2_1 U23169 ( .ip1(\x[64][10] ), .ip2(n23980), .op(n19150) );
  nand2_1 U23170 ( .ip1(n19151), .ip2(n19150), .op(n19154) );
  inv_1 U23171 ( .ip(n19152), .op(n19153) );
  nand2_1 U23172 ( .ip1(n19154), .ip2(n19153), .op(n19157) );
  nand2_1 U23173 ( .ip1(\x[64][13] ), .ip2(n24081), .op(n19156) );
  nand2_1 U23174 ( .ip1(\x[64][14] ), .ip2(n24327), .op(n19155) );
  nand4_1 U23175 ( .ip1(n19158), .ip2(n19157), .ip3(n19156), .ip4(n19155), 
        .op(n19160) );
  or2_1 U23176 ( .ip1(n19160), .ip2(n19159), .op(n19161) );
  nand2_1 U23177 ( .ip1(n19162), .ip2(n19161), .op(n19277) );
  inv_1 U23178 ( .ip(n19163), .op(n19164) );
  nand2_1 U23179 ( .ip1(n19165), .ip2(n19164), .op(n19167) );
  nand2_1 U23180 ( .ip1(n19167), .ip2(n19166), .op(n19169) );
  nand2_1 U23181 ( .ip1(n19169), .ip2(n19168), .op(n19176) );
  or3_1 U23182 ( .ip1(n19171), .ip2(n19170), .ip3(n17845), .op(n19175) );
  or2_1 U23183 ( .ip1(n19173), .ip2(n19172), .op(n19174) );
  nand4_1 U23184 ( .ip1(n19277), .ip2(n19176), .ip3(n19175), .ip4(n19174), 
        .op(n24674) );
  nand2_1 U23185 ( .ip1(n24672), .ip2(n24674), .op(n24687) );
  nand2_1 U23186 ( .ip1(\x[62][15] ), .ip2(n24186), .op(n19257) );
  and2_1 U23187 ( .ip1(n23895), .ip2(\x[62][13] ), .op(n19177) );
  nor2_1 U23188 ( .ip1(\x[62][15] ), .ip2(n23143), .op(n19301) );
  not_ab_or_c_or_d U23189 ( .ip1(\x[62][14] ), .ip2(n23938), .ip3(n19177), 
        .ip4(n19301), .op(n19299) );
  nand2_1 U23190 ( .ip1(\x[62][12] ), .ip2(n24233), .op(n19296) );
  nand2_1 U23191 ( .ip1(n19299), .ip2(n19296), .op(n19256) );
  and2_1 U23192 ( .ip1(n24451), .ip2(\x[63][10] ), .op(n19179) );
  and2_1 U23193 ( .ip1(n24239), .ip2(\x[63][11] ), .op(n19178) );
  not_ab_or_c_or_d U23194 ( .ip1(\x[63][9] ), .ip2(n23981), .ip3(n19179), 
        .ip4(n19178), .op(n19261) );
  nor2_1 U23195 ( .ip1(n24371), .ip2(\x[63][11] ), .op(n19181) );
  not_ab_or_c_or_d U23196 ( .ip1(\x[63][11] ), .ip2(n24136), .ip3(\x[63][10] ), 
        .ip4(n20880), .op(n19180) );
  or2_1 U23197 ( .ip1(n19181), .ip2(n19180), .op(n19270) );
  or2_1 U23198 ( .ip1(n19261), .ip2(n19270), .op(n19207) );
  nor2_1 U23199 ( .ip1(\x[63][9] ), .ip2(n23981), .op(n19260) );
  or2_1 U23200 ( .ip1(n23779), .ip2(n19260), .op(n19184) );
  inv_1 U23201 ( .ip(\x[63][8] ), .op(n19182) );
  or2_1 U23202 ( .ip1(n19182), .ip2(n19260), .op(n19183) );
  nand2_1 U23203 ( .ip1(n19184), .ip2(n19183), .op(n19265) );
  nor2_1 U23204 ( .ip1(n24142), .ip2(\x[63][7] ), .op(n19202) );
  inv_1 U23205 ( .ip(\x[63][5] ), .op(n19198) );
  nor2_1 U23206 ( .ip1(n22833), .ip2(n19198), .op(n19195) );
  inv_1 U23207 ( .ip(\x[63][3] ), .op(n19193) );
  inv_1 U23208 ( .ip(n24251), .op(n24476) );
  and2_1 U23209 ( .ip1(n24335), .ip2(\x[63][2] ), .op(n19190) );
  inv_1 U23210 ( .ip(sig_in[1]), .op(n21685) );
  nand2_1 U23211 ( .ip1(\x[63][1] ), .ip2(n21685), .op(n19188) );
  nand2_1 U23212 ( .ip1(\x[63][0] ), .ip2(n24143), .op(n19187) );
  nor2_1 U23213 ( .ip1(\x[63][2] ), .ip2(n24463), .op(n19186) );
  nor2_1 U23214 ( .ip1(\x[63][1] ), .ip2(n21685), .op(n19185) );
  not_ab_or_c_or_d U23215 ( .ip1(n19188), .ip2(n19187), .ip3(n19186), .ip4(
        n19185), .op(n19189) );
  not_ab_or_c_or_d U23216 ( .ip1(\x[63][3] ), .ip2(n24476), .ip3(n19190), 
        .ip4(n19189), .op(n19192) );
  nor2_1 U23217 ( .ip1(\x[63][4] ), .ip2(n23721), .op(n19191) );
  not_ab_or_c_or_d U23218 ( .ip1(n23251), .ip2(n19193), .ip3(n19192), .ip4(
        n19191), .op(n19194) );
  not_ab_or_c_or_d U23219 ( .ip1(\x[63][4] ), .ip2(n23860), .ip3(n19195), 
        .ip4(n19194), .op(n19197) );
  nor2_1 U23220 ( .ip1(\x[63][6] ), .ip2(n24355), .op(n19196) );
  not_ab_or_c_or_d U23221 ( .ip1(n22833), .ip2(n19198), .ip3(n19197), .ip4(
        n19196), .op(n19200) );
  and2_1 U23222 ( .ip1(n23509), .ip2(\x[63][6] ), .op(n19199) );
  not_ab_or_c_or_d U23223 ( .ip1(\x[63][7] ), .ip2(n24142), .ip3(n19200), 
        .ip4(n19199), .op(n19201) );
  nor2_1 U23224 ( .ip1(n19202), .ip2(n19201), .op(n19264) );
  inv_1 U23225 ( .ip(n19264), .op(n19203) );
  nand2_1 U23226 ( .ip1(\x[63][8] ), .ip2(n23804), .op(n19259) );
  nand2_1 U23227 ( .ip1(n19203), .ip2(n19259), .op(n19204) );
  nand2_1 U23228 ( .ip1(n19265), .ip2(n19204), .op(n19205) );
  or2_1 U23229 ( .ip1(n19205), .ip2(n19270), .op(n19206) );
  nand2_1 U23230 ( .ip1(n19207), .ip2(n19206), .op(n19210) );
  and2_1 U23231 ( .ip1(n23895), .ip2(\x[63][13] ), .op(n19208) );
  nor2_1 U23232 ( .ip1(\x[63][15] ), .ip2(n23143), .op(n19216) );
  not_ab_or_c_or_d U23233 ( .ip1(\x[63][14] ), .ip2(n24327), .ip3(n19208), 
        .ip4(n19216), .op(n19253) );
  nand2_1 U23234 ( .ip1(\x[63][12] ), .ip2(n24449), .op(n19209) );
  nand2_1 U23235 ( .ip1(n19253), .ip2(n19209), .op(n19271) );
  nor2_1 U23236 ( .ip1(n19210), .ip2(n19271), .op(n19255) );
  nor2_1 U23237 ( .ip1(\x[63][13] ), .ip2(n24081), .op(n19212) );
  nor2_1 U23238 ( .ip1(\x[63][12] ), .ip2(n24449), .op(n19211) );
  or2_1 U23239 ( .ip1(n19212), .ip2(n19211), .op(n19267) );
  and2_1 U23240 ( .ip1(n24186), .ip2(\x[63][15] ), .op(n19272) );
  or2_1 U23241 ( .ip1(sig_in[14]), .ip2(n19272), .op(n19215) );
  inv_1 U23242 ( .ip(\x[63][14] ), .op(n19213) );
  or2_1 U23243 ( .ip1(n19213), .ip2(n19272), .op(n19214) );
  nand2_1 U23244 ( .ip1(n19215), .ip2(n19214), .op(n19266) );
  nor2_1 U23245 ( .ip1(n19216), .ip2(n19266), .op(n19252) );
  inv_1 U23246 ( .ip(\x[62][11] ), .op(n19243) );
  and2_1 U23247 ( .ip1(n24451), .ip2(\x[62][10] ), .op(n19240) );
  nor2_1 U23248 ( .ip1(\x[62][7] ), .ip2(n24142), .op(n19231) );
  inv_1 U23249 ( .ip(\x[62][6] ), .op(n19217) );
  nor3_1 U23250 ( .ip1(sig_in[6]), .ip2(n19231), .ip3(n19217), .op(n19234) );
  and2_1 U23251 ( .ip1(n23283), .ip2(\x[62][5] ), .op(n19228) );
  inv_1 U23252 ( .ip(\x[62][3] ), .op(n19226) );
  and2_1 U23253 ( .ip1(n24335), .ip2(\x[62][2] ), .op(n19223) );
  inv_1 U23254 ( .ip(sig_in[0]), .op(n24143) );
  nand3_1 U23255 ( .ip1(\x[62][0] ), .ip2(\x[62][1] ), .ip3(n24143), .op(
        n19221) );
  nor2_1 U23256 ( .ip1(\x[62][2] ), .ip2(n23717), .op(n19220) );
  and2_1 U23257 ( .ip1(n24143), .ip2(\x[62][0] ), .op(n19218) );
  nor2_1 U23258 ( .ip1(n19218), .ip2(\x[62][1] ), .op(n19219) );
  not_ab_or_c_or_d U23259 ( .ip1(n24464), .ip2(n19221), .ip3(n19220), .ip4(
        n19219), .op(n19222) );
  not_ab_or_c_or_d U23260 ( .ip1(\x[62][3] ), .ip2(n24476), .ip3(n19223), 
        .ip4(n19222), .op(n19225) );
  nor2_1 U23261 ( .ip1(\x[62][4] ), .ip2(n24256), .op(n19224) );
  not_ab_or_c_or_d U23262 ( .ip1(n24251), .ip2(n19226), .ip3(n19225), .ip4(
        n19224), .op(n19227) );
  not_ab_or_c_or_d U23263 ( .ip1(\x[62][4] ), .ip2(n23860), .ip3(n19228), 
        .ip4(n19227), .op(n19232) );
  nor2_1 U23264 ( .ip1(\x[62][5] ), .ip2(n23283), .op(n19230) );
  nor2_1 U23265 ( .ip1(\x[62][6] ), .ip2(n23509), .op(n19229) );
  nor4_1 U23266 ( .ip1(n19232), .ip2(n19231), .ip3(n19230), .ip4(n19229), .op(
        n19233) );
  not_ab_or_c_or_d U23267 ( .ip1(\x[62][7] ), .ip2(n24492), .ip3(n19234), 
        .ip4(n19233), .op(n19238) );
  nand2_1 U23268 ( .ip1(\x[62][8] ), .ip2(n24491), .op(n19237) );
  nor2_1 U23269 ( .ip1(\x[62][9] ), .ip2(n24164), .op(n19236) );
  nor2_1 U23270 ( .ip1(\x[62][8] ), .ip2(n23971), .op(n19235) );
  not_ab_or_c_or_d U23271 ( .ip1(n19238), .ip2(n19237), .ip3(n19236), .ip4(
        n19235), .op(n19239) );
  not_ab_or_c_or_d U23272 ( .ip1(\x[62][9] ), .ip2(n23981), .ip3(n19240), 
        .ip4(n19239), .op(n19242) );
  nor2_1 U23273 ( .ip1(\x[62][10] ), .ip2(n20880), .op(n19241) );
  not_ab_or_c_or_d U23274 ( .ip1(sig_in[11]), .ip2(n19243), .ip3(n19242), 
        .ip4(n19241), .op(n19244) );
  or2_1 U23275 ( .ip1(\x[62][11] ), .ip2(n19244), .op(n19246) );
  or2_1 U23276 ( .ip1(n24136), .ip2(n19244), .op(n19245) );
  nand2_1 U23277 ( .ip1(n19246), .ip2(n19245), .op(n19295) );
  nor2_1 U23278 ( .ip1(\x[62][13] ), .ip2(n23895), .op(n19248) );
  nor2_1 U23279 ( .ip1(\x[62][12] ), .ip2(n24449), .op(n19247) );
  nor2_1 U23280 ( .ip1(n19248), .ip2(n19247), .op(n19297) );
  inv_1 U23281 ( .ip(n19297), .op(n19250) );
  or2_1 U23282 ( .ip1(n24185), .ip2(\x[62][14] ), .op(n19249) );
  nand2_1 U23283 ( .ip1(n19257), .ip2(n19249), .op(n19303) );
  nor3_1 U23284 ( .ip1(n19295), .ip2(n19250), .ip3(n19303), .op(n19251) );
  ab_or_c_or_d U23285 ( .ip1(n19253), .ip2(n19267), .ip3(n19252), .ip4(n19251), 
        .op(n19254) );
  ab_or_c_or_d U23286 ( .ip1(n19257), .ip2(n19256), .ip3(n19255), .ip4(n19254), 
        .op(n24686) );
  nand3_1 U23287 ( .ip1(\x[64][12] ), .ip2(n19258), .ip3(n24450), .op(n19276)
         );
  nor2_1 U23288 ( .ip1(n19260), .ip2(n19259), .op(n19263) );
  inv_1 U23289 ( .ip(n19261), .op(n19262) );
  not_ab_or_c_or_d U23290 ( .ip1(n19265), .ip2(n19264), .ip3(n19263), .ip4(
        n19262), .op(n19269) );
  inv_1 U23291 ( .ip(n19266), .op(n19268) );
  nor4_1 U23292 ( .ip1(n19270), .ip2(n19269), .ip3(n19268), .ip4(n19267), .op(
        n19275) );
  inv_1 U23293 ( .ip(n19271), .op(n19273) );
  nor2_1 U23294 ( .ip1(n19273), .ip2(n19272), .op(n19274) );
  ab_or_c_or_d U23295 ( .ip1(n19277), .ip2(n19276), .ip3(n19275), .ip4(n19274), 
        .op(n24678) );
  nand2_1 U23296 ( .ip1(n24686), .ip2(n24678), .op(n19278) );
  nor2_1 U23297 ( .ip1(n24687), .ip2(n19278), .op(n24688) );
  inv_1 U23298 ( .ip(n19279), .op(n19287) );
  not_ab_or_c_or_d U23299 ( .ip1(n19283), .ip2(n19282), .ip3(n19281), .ip4(
        n19280), .op(n19285) );
  not_ab_or_c_or_d U23300 ( .ip1(n19287), .ip2(n19286), .ip3(n19285), .ip4(
        n19284), .op(n19292) );
  nand3_1 U23301 ( .ip1(n19290), .ip2(n19289), .ip3(n19288), .op(n19291) );
  nand2_1 U23302 ( .ip1(n19292), .ip2(n19291), .op(n19293) );
  nand2_1 U23303 ( .ip1(n19294), .ip2(n19293), .op(n19306) );
  nand2_1 U23304 ( .ip1(n19296), .ip2(n19295), .op(n19298) );
  nand2_1 U23305 ( .ip1(n19298), .ip2(n19297), .op(n19300) );
  nand2_1 U23306 ( .ip1(n19300), .ip2(n19299), .op(n19305) );
  inv_1 U23307 ( .ip(n19301), .op(n19302) );
  nand2_1 U23308 ( .ip1(n19303), .ip2(n19302), .op(n19304) );
  nand3_1 U23309 ( .ip1(n19306), .ip2(n19305), .ip3(n19304), .op(n24690) );
  nand2_1 U23310 ( .ip1(n24688), .ip2(n24690), .op(n24692) );
  nor2_1 U23311 ( .ip1(n24691), .ip2(n24692), .op(n24675) );
  or2_1 U23312 ( .ip1(n19308), .ip2(n19307), .op(n19318) );
  inv_1 U23313 ( .ip(n19309), .op(n19310) );
  nand2_1 U23314 ( .ip1(n19311), .ip2(n19310), .op(n19313) );
  nand2_1 U23315 ( .ip1(n19313), .ip2(n19312), .op(n19315) );
  nand2_1 U23316 ( .ip1(n19315), .ip2(n19314), .op(n19317) );
  nand3_1 U23317 ( .ip1(n19318), .ip2(n19317), .ip3(n19316), .op(n24677) );
  nand2_1 U23318 ( .ip1(n24675), .ip2(n24677), .op(n24652) );
  or2_1 U23319 ( .ip1(n24651), .ip2(n24652), .op(n24684) );
  nor2_1 U23320 ( .ip1(n24683), .ip2(n24684), .op(n26760) );
  or2_1 U23321 ( .ip1(n19320), .ip2(n19319), .op(n19323) );
  nand3_1 U23322 ( .ip1(n19323), .ip2(n19322), .ip3(n19321), .op(n19377) );
  and2_1 U23323 ( .ip1(n24186), .ip2(\x[44][15] ), .op(n20046) );
  or2_1 U23324 ( .ip1(sig_in[14]), .ip2(n20046), .op(n19326) );
  inv_1 U23325 ( .ip(\x[44][14] ), .op(n19324) );
  or2_1 U23326 ( .ip1(n19324), .ip2(n20046), .op(n19325) );
  nand2_1 U23327 ( .ip1(n19326), .ip2(n19325), .op(n20035) );
  nor2_1 U23328 ( .ip1(\x[44][15] ), .ip2(n24090), .op(n19369) );
  nor2_1 U23329 ( .ip1(n20035), .ip2(n19369), .op(n19376) );
  inv_1 U23330 ( .ip(\x[44][11] ), .op(n19357) );
  nand2_1 U23331 ( .ip1(\x[44][9] ), .ip2(n24455), .op(n19329) );
  nand2_1 U23332 ( .ip1(\x[44][8] ), .ip2(n24100), .op(n19327) );
  nor2_1 U23333 ( .ip1(\x[44][9] ), .ip2(n24043), .op(n19351) );
  or2_1 U23334 ( .ip1(n19327), .ip2(n19351), .op(n19328) );
  nand2_1 U23335 ( .ip1(n19329), .ip2(n19328), .op(n19354) );
  nor2_1 U23336 ( .ip1(\x[44][7] ), .ip2(n24492), .op(n19352) );
  nor2_1 U23337 ( .ip1(\x[44][8] ), .ip2(n24358), .op(n19350) );
  and2_1 U23338 ( .ip1(n24461), .ip2(\x[44][7] ), .op(n19346) );
  nor3_1 U23339 ( .ip1(n24045), .ip2(\x[44][6] ), .ip3(n19346), .op(n19348) );
  inv_1 U23340 ( .ip(\x[44][3] ), .op(n19336) );
  nor2_1 U23341 ( .ip1(n19336), .ip2(sig_in[3]), .op(n19338) );
  inv_1 U23342 ( .ip(\x[44][1] ), .op(n19331) );
  nor2_1 U23343 ( .ip1(n22513), .ip2(n19331), .op(n19333) );
  inv_1 U23344 ( .ip(\x[44][0] ), .op(n19330) );
  not_ab_or_c_or_d U23345 ( .ip1(n24464), .ip2(n19331), .ip3(sig_in[0]), .ip4(
        n19330), .op(n19332) );
  not_ab_or_c_or_d U23346 ( .ip1(\x[44][2] ), .ip2(n24107), .ip3(n19333), 
        .ip4(n19332), .op(n19335) );
  nor2_1 U23347 ( .ip1(\x[44][2] ), .ip2(n23717), .op(n19334) );
  not_ab_or_c_or_d U23348 ( .ip1(sig_in[3]), .ip2(n19336), .ip3(n19335), .ip4(
        n19334), .op(n19337) );
  or2_1 U23349 ( .ip1(n19338), .ip2(n19337), .op(n19339) );
  nand2_1 U23350 ( .ip1(\x[44][4] ), .ip2(n19339), .op(n19342) );
  nor2_1 U23351 ( .ip1(\x[44][5] ), .ip2(n23600), .op(n19341) );
  nor2_1 U23352 ( .ip1(\x[44][4] ), .ip2(n19339), .op(n19340) );
  ab_or_c_or_d U23353 ( .ip1(sig_in[4]), .ip2(n19342), .ip3(n19341), .ip4(
        n19340), .op(n19344) );
  nand2_1 U23354 ( .ip1(\x[44][5] ), .ip2(n24119), .op(n19343) );
  nand2_1 U23355 ( .ip1(n19344), .ip2(n19343), .op(n19345) );
  not_ab_or_c_or_d U23356 ( .ip1(\x[44][6] ), .ip2(n24355), .ip3(n19346), 
        .ip4(n19345), .op(n19347) );
  or2_1 U23357 ( .ip1(n19348), .ip2(n19347), .op(n19349) );
  nor4_1 U23358 ( .ip1(n19352), .ip2(n19351), .ip3(n19350), .ip4(n19349), .op(
        n19353) );
  not_ab_or_c_or_d U23359 ( .ip1(\x[44][10] ), .ip2(n23980), .ip3(n19354), 
        .ip4(n19353), .op(n19356) );
  buf_1 U23360 ( .ip(n24370), .op(n24457) );
  nor2_1 U23361 ( .ip1(\x[44][10] ), .ip2(n24457), .op(n19355) );
  not_ab_or_c_or_d U23362 ( .ip1(sig_in[11]), .ip2(n19357), .ip3(n19356), 
        .ip4(n19355), .op(n19358) );
  or2_1 U23363 ( .ip1(\x[44][11] ), .ip2(n19358), .op(n19360) );
  or2_1 U23364 ( .ip1(n24136), .ip2(n19358), .op(n19359) );
  nand2_1 U23365 ( .ip1(n19360), .ip2(n19359), .op(n20040) );
  and2_1 U23366 ( .ip1(n24332), .ip2(\x[44][13] ), .op(n19361) );
  or2_1 U23367 ( .ip1(\x[44][12] ), .ip2(n19361), .op(n19363) );
  or2_1 U23368 ( .ip1(n24233), .ip2(n19361), .op(n19362) );
  nand2_1 U23369 ( .ip1(n19363), .ip2(n19362), .op(n20036) );
  nand2_1 U23370 ( .ip1(n20040), .ip2(n20036), .op(n19368) );
  nor2_1 U23371 ( .ip1(\x[44][13] ), .ip2(n24332), .op(n19364) );
  or2_1 U23372 ( .ip1(sig_in[12]), .ip2(n19364), .op(n19367) );
  inv_1 U23373 ( .ip(\x[44][12] ), .op(n19365) );
  or2_1 U23374 ( .ip1(n19365), .ip2(n19364), .op(n19366) );
  nand2_1 U23375 ( .ip1(n19367), .ip2(n19366), .op(n20037) );
  nand2_1 U23376 ( .ip1(n19368), .ip2(n20037), .op(n19372) );
  or2_1 U23377 ( .ip1(\x[44][14] ), .ip2(n19369), .op(n19371) );
  or2_1 U23378 ( .ip1(n24185), .ip2(n19369), .op(n19370) );
  nand2_1 U23379 ( .ip1(n19371), .ip2(n19370), .op(n20045) );
  nand2_1 U23380 ( .ip1(n19372), .ip2(n20045), .op(n19374) );
  nand2_1 U23381 ( .ip1(n19374), .ip2(n19373), .op(n19375) );
  not_ab_or_c_or_d U23382 ( .ip1(n19378), .ip2(n19377), .ip3(n19376), .ip4(
        n19375), .op(n24835) );
  nand2_1 U23383 ( .ip1(\x[46][15] ), .ip2(n24180), .op(n19474) );
  or2_1 U23384 ( .ip1(n24384), .ip2(\x[46][15] ), .op(n20026) );
  nand2_1 U23385 ( .ip1(\x[46][14] ), .ip2(n24327), .op(n19379) );
  nand2_1 U23386 ( .ip1(n20026), .ip2(n19379), .op(n20029) );
  nor2_1 U23387 ( .ip1(\x[47][15] ), .ip2(n23143), .op(n19429) );
  nor2_1 U23388 ( .ip1(\x[47][14] ), .ip2(n24230), .op(n19380) );
  or2_1 U23389 ( .ip1(\x[47][15] ), .ip2(n19380), .op(n19382) );
  or2_1 U23390 ( .ip1(n24384), .ip2(n19380), .op(n19381) );
  nand2_1 U23391 ( .ip1(n19382), .ip2(n19381), .op(n19977) );
  nor2_1 U23392 ( .ip1(n19429), .ip2(n19977), .op(n19966) );
  or2_1 U23393 ( .ip1(n24382), .ip2(\x[46][14] ), .op(n19383) );
  nand2_1 U23394 ( .ip1(n19474), .ip2(n19383), .op(n20027) );
  nand2_1 U23395 ( .ip1(\x[46][13] ), .ip2(n24081), .op(n19385) );
  nand2_1 U23396 ( .ip1(\x[46][12] ), .ip2(n24450), .op(n19384) );
  nand2_1 U23397 ( .ip1(n19385), .ip2(n19384), .op(n20028) );
  inv_1 U23398 ( .ip(\x[46][12] ), .op(n19423) );
  nor2_1 U23399 ( .ip1(\x[46][9] ), .ip2(n24269), .op(n19410) );
  inv_1 U23400 ( .ip(\x[46][8] ), .op(n19386) );
  nor3_1 U23401 ( .ip1(sig_in[8]), .ip2(n19410), .ip3(n19386), .op(n19413) );
  and2_1 U23402 ( .ip1(n24461), .ip2(\x[46][7] ), .op(n19407) );
  inv_1 U23403 ( .ip(\x[46][5] ), .op(n19405) );
  nor2_1 U23404 ( .ip1(n22833), .ip2(n19405), .op(n19402) );
  inv_1 U23405 ( .ip(\x[46][3] ), .op(n19393) );
  inv_1 U23406 ( .ip(\x[46][1] ), .op(n19388) );
  nor2_1 U23407 ( .ip1(n22513), .ip2(n19388), .op(n19390) );
  buf_1 U23408 ( .ip(sig_in[0]), .op(n23195) );
  inv_1 U23409 ( .ip(\x[46][0] ), .op(n19387) );
  not_ab_or_c_or_d U23410 ( .ip1(n24467), .ip2(n19388), .ip3(n23195), .ip4(
        n19387), .op(n19389) );
  not_ab_or_c_or_d U23411 ( .ip1(\x[46][2] ), .ip2(n24107), .ip3(n19390), 
        .ip4(n19389), .op(n19392) );
  nor2_1 U23412 ( .ip1(\x[46][2] ), .ip2(n23717), .op(n19391) );
  not_ab_or_c_or_d U23413 ( .ip1(sig_in[3]), .ip2(n19393), .ip3(n19392), .ip4(
        n19391), .op(n19394) );
  or2_1 U23414 ( .ip1(\x[46][3] ), .ip2(n19394), .op(n19396) );
  or2_1 U23415 ( .ip1(n24476), .ip2(n19394), .op(n19395) );
  nand2_1 U23416 ( .ip1(n19396), .ip2(n19395), .op(n19397) );
  or2_1 U23417 ( .ip1(sig_in[4]), .ip2(n19397), .op(n19400) );
  inv_1 U23418 ( .ip(\x[46][4] ), .op(n19398) );
  or2_1 U23419 ( .ip1(n19398), .ip2(n19397), .op(n19399) );
  nand2_1 U23420 ( .ip1(n19400), .ip2(n19399), .op(n19401) );
  not_ab_or_c_or_d U23421 ( .ip1(\x[46][4] ), .ip2(n23860), .ip3(n19402), 
        .ip4(n19401), .op(n19404) );
  nor2_1 U23422 ( .ip1(\x[46][6] ), .ip2(n23509), .op(n19403) );
  not_ab_or_c_or_d U23423 ( .ip1(n22833), .ip2(n19405), .ip3(n19404), .ip4(
        n19403), .op(n19406) );
  not_ab_or_c_or_d U23424 ( .ip1(\x[46][6] ), .ip2(n24355), .ip3(n19407), 
        .ip4(n19406), .op(n19411) );
  nor2_1 U23425 ( .ip1(\x[46][8] ), .ip2(n23971), .op(n19409) );
  nor2_1 U23426 ( .ip1(\x[46][7] ), .ip2(n24044), .op(n19408) );
  nor4_1 U23427 ( .ip1(n19411), .ip2(n19410), .ip3(n19409), .ip4(n19408), .op(
        n19412) );
  not_ab_or_c_or_d U23428 ( .ip1(\x[46][10] ), .ip2(n24370), .ip3(n19413), 
        .ip4(n19412), .op(n19417) );
  nand2_1 U23429 ( .ip1(\x[46][9] ), .ip2(n23981), .op(n19416) );
  nor2_1 U23430 ( .ip1(\x[46][11] ), .ip2(n24371), .op(n19415) );
  nor2_1 U23431 ( .ip1(\x[46][10] ), .ip2(n20880), .op(n19414) );
  not_ab_or_c_or_d U23432 ( .ip1(n19417), .ip2(n19416), .ip3(n19415), .ip4(
        n19414), .op(n19418) );
  or2_1 U23433 ( .ip1(\x[46][11] ), .ip2(n19418), .op(n19420) );
  or2_1 U23434 ( .ip1(n24136), .ip2(n19418), .op(n19419) );
  nand2_1 U23435 ( .ip1(n19420), .ip2(n19419), .op(n19422) );
  nor2_1 U23436 ( .ip1(\x[46][13] ), .ip2(n24235), .op(n19421) );
  not_ab_or_c_or_d U23437 ( .ip1(sig_in[12]), .ip2(n19423), .ip3(n19422), 
        .ip4(n19421), .op(n20030) );
  nor2_1 U23438 ( .ip1(n20028), .ip2(n20030), .op(n19424) );
  nor2_1 U23439 ( .ip1(n20027), .ip2(n19424), .op(n19434) );
  nor2_1 U23440 ( .ip1(\x[47][13] ), .ip2(n24137), .op(n19425) );
  or2_1 U23441 ( .ip1(sig_in[12]), .ip2(n19425), .op(n19428) );
  inv_1 U23442 ( .ip(\x[47][12] ), .op(n19426) );
  or2_1 U23443 ( .ip1(n19426), .ip2(n19425), .op(n19427) );
  nand2_1 U23444 ( .ip1(n19428), .ip2(n19427), .op(n19975) );
  nand2_1 U23445 ( .ip1(n24185), .ip2(\x[47][14] ), .op(n19432) );
  inv_1 U23446 ( .ip(n19429), .op(n19431) );
  nand2_1 U23447 ( .ip1(\x[47][13] ), .ip2(n24235), .op(n19430) );
  nand3_1 U23448 ( .ip1(n19432), .ip2(n19431), .ip3(n19430), .op(n19435) );
  nor2_1 U23449 ( .ip1(n19975), .ip2(n19435), .op(n19433) );
  nor2_1 U23450 ( .ip1(n19434), .ip2(n19433), .op(n19472) );
  or2_1 U23451 ( .ip1(\x[47][12] ), .ip2(n19435), .op(n19437) );
  or2_1 U23452 ( .ip1(n24233), .ip2(n19435), .op(n19436) );
  nand2_1 U23453 ( .ip1(n19437), .ip2(n19436), .op(n19967) );
  and2_1 U23454 ( .ip1(n24371), .ip2(\x[47][11] ), .op(n19470) );
  nor2_1 U23455 ( .ip1(\x[47][10] ), .ip2(n20880), .op(n19468) );
  and2_1 U23456 ( .ip1(n23146), .ip2(\x[47][10] ), .op(n19465) );
  inv_1 U23457 ( .ip(\x[47][9] ), .op(n19463) );
  nor2_1 U23458 ( .ip1(\x[47][8] ), .ip2(n23971), .op(n19462) );
  inv_1 U23459 ( .ip(sig_in[8]), .op(n23804) );
  and2_1 U23460 ( .ip1(n23804), .ip2(\x[47][8] ), .op(n19460) );
  inv_1 U23461 ( .ip(\x[47][5] ), .op(n19451) );
  nor2_1 U23462 ( .ip1(n22833), .ip2(n19451), .op(n19448) );
  inv_1 U23463 ( .ip(\x[47][3] ), .op(n19446) );
  buf_1 U23464 ( .ip(n24107), .op(n23659) );
  and2_1 U23465 ( .ip1(n23659), .ip2(\x[47][2] ), .op(n19443) );
  nand2_1 U23466 ( .ip1(\x[47][1] ), .ip2(n21685), .op(n19441) );
  nand2_1 U23467 ( .ip1(\x[47][0] ), .ip2(n24143), .op(n19440) );
  nor2_1 U23468 ( .ip1(\x[47][2] ), .ip2(n24463), .op(n19439) );
  nor2_1 U23469 ( .ip1(\x[47][1] ), .ip2(n21685), .op(n19438) );
  not_ab_or_c_or_d U23470 ( .ip1(n19441), .ip2(n19440), .ip3(n19439), .ip4(
        n19438), .op(n19442) );
  not_ab_or_c_or_d U23471 ( .ip1(\x[47][3] ), .ip2(n22525), .ip3(n19443), 
        .ip4(n19442), .op(n19445) );
  nor2_1 U23472 ( .ip1(\x[47][4] ), .ip2(n23721), .op(n19444) );
  not_ab_or_c_or_d U23473 ( .ip1(sig_in[3]), .ip2(n19446), .ip3(n19445), .ip4(
        n19444), .op(n19447) );
  not_ab_or_c_or_d U23474 ( .ip1(\x[47][4] ), .ip2(n23860), .ip3(n19448), 
        .ip4(n19447), .op(n19450) );
  nor2_1 U23475 ( .ip1(\x[47][6] ), .ip2(n23509), .op(n19449) );
  not_ab_or_c_or_d U23476 ( .ip1(n22833), .ip2(n19451), .ip3(n19450), .ip4(
        n19449), .op(n19452) );
  or2_1 U23477 ( .ip1(\x[47][6] ), .ip2(n19452), .op(n19454) );
  or2_1 U23478 ( .ip1(n24045), .ip2(n19452), .op(n19453) );
  nand2_1 U23479 ( .ip1(n19454), .ip2(n19453), .op(n19455) );
  or2_1 U23480 ( .ip1(sig_in[7]), .ip2(n19455), .op(n19458) );
  inv_1 U23481 ( .ip(\x[47][7] ), .op(n19456) );
  or2_1 U23482 ( .ip1(n19456), .ip2(n19455), .op(n19457) );
  nand2_1 U23483 ( .ip1(n19458), .ip2(n19457), .op(n19459) );
  not_ab_or_c_or_d U23484 ( .ip1(\x[47][7] ), .ip2(n24492), .ip3(n19460), 
        .ip4(n19459), .op(n19461) );
  not_ab_or_c_or_d U23485 ( .ip1(n21171), .ip2(n19463), .ip3(n19462), .ip4(
        n19461), .op(n19464) );
  not_ab_or_c_or_d U23486 ( .ip1(\x[47][9] ), .ip2(n23981), .ip3(n19465), 
        .ip4(n19464), .op(n19467) );
  nor2_1 U23487 ( .ip1(\x[47][11] ), .ip2(n24371), .op(n19466) );
  nor3_1 U23488 ( .ip1(n19468), .ip2(n19467), .ip3(n19466), .op(n19469) );
  nor2_1 U23489 ( .ip1(n19470), .ip2(n19469), .op(n19974) );
  nand2_1 U23490 ( .ip1(n19967), .ip2(n19974), .op(n19471) );
  nand2_1 U23491 ( .ip1(n19472), .ip2(n19471), .op(n19473) );
  not_ab_or_c_or_d U23492 ( .ip1(n19474), .ip2(n20029), .ip3(n19966), .ip4(
        n19473), .op(n24800) );
  and2_1 U23493 ( .ip1(n24332), .ip2(\x[49][13] ), .op(n19475) );
  nor2_1 U23494 ( .ip1(\x[49][15] ), .ip2(n23143), .op(n19482) );
  not_ab_or_c_or_d U23495 ( .ip1(\x[49][14] ), .ip2(n24230), .ip3(n19475), 
        .ip4(n19482), .op(n19575) );
  nor2_1 U23496 ( .ip1(\x[49][13] ), .ip2(n24376), .op(n19477) );
  nor2_1 U23497 ( .ip1(\x[49][12] ), .ip2(n24449), .op(n19476) );
  or2_1 U23498 ( .ip1(n19477), .ip2(n19476), .op(n19636) );
  nand2_1 U23499 ( .ip1(n24384), .ip2(\x[49][15] ), .op(n19640) );
  inv_1 U23500 ( .ip(n19640), .op(n19478) );
  or2_1 U23501 ( .ip1(sig_in[14]), .ip2(n19478), .op(n19481) );
  inv_1 U23502 ( .ip(\x[49][14] ), .op(n19479) );
  or2_1 U23503 ( .ip1(n19479), .ip2(n19478), .op(n19480) );
  nand2_1 U23504 ( .ip1(n19481), .ip2(n19480), .op(n19634) );
  nor2_1 U23505 ( .ip1(n19482), .ip2(n19634), .op(n19574) );
  and2_1 U23506 ( .ip1(\x[49][11] ), .ip2(n24371), .op(n19513) );
  nor2_1 U23507 ( .ip1(\x[49][11] ), .ip2(n24239), .op(n19484) );
  nor2_1 U23508 ( .ip1(\x[49][10] ), .ip2(n20880), .op(n19483) );
  nor2_1 U23509 ( .ip1(n19484), .ip2(n19483), .op(n19633) );
  or2_1 U23510 ( .ip1(n19513), .ip2(n19633), .op(n19630) );
  nor2_1 U23511 ( .ip1(n24142), .ip2(\x[49][7] ), .op(n19507) );
  inv_1 U23512 ( .ip(\x[49][5] ), .op(n19503) );
  inv_1 U23513 ( .ip(\x[49][4] ), .op(n19495) );
  nor2_1 U23514 ( .ip1(n24462), .ip2(n19495), .op(n19493) );
  inv_1 U23515 ( .ip(\x[49][3] ), .op(n19491) );
  inv_1 U23516 ( .ip(\x[49][1] ), .op(n19486) );
  nor2_1 U23517 ( .ip1(n22513), .ip2(n19486), .op(n19488) );
  inv_1 U23518 ( .ip(\x[49][0] ), .op(n19485) );
  not_ab_or_c_or_d U23519 ( .ip1(n24464), .ip2(n19486), .ip3(n23195), .ip4(
        n19485), .op(n19487) );
  not_ab_or_c_or_d U23520 ( .ip1(\x[49][2] ), .ip2(n24470), .ip3(n19488), 
        .ip4(n19487), .op(n19490) );
  nor2_1 U23521 ( .ip1(\x[49][2] ), .ip2(n23717), .op(n19489) );
  not_ab_or_c_or_d U23522 ( .ip1(sig_in[3]), .ip2(n19491), .ip3(n19490), .ip4(
        n19489), .op(n19492) );
  not_ab_or_c_or_d U23523 ( .ip1(\x[49][3] ), .ip2(n24476), .ip3(n19493), 
        .ip4(n19492), .op(n19494) );
  or2_1 U23524 ( .ip1(sig_in[4]), .ip2(n19494), .op(n19497) );
  or2_1 U23525 ( .ip1(n19495), .ip2(n19494), .op(n19496) );
  nand2_1 U23526 ( .ip1(n19497), .ip2(n19496), .op(n19498) );
  or2_1 U23527 ( .ip1(\x[49][5] ), .ip2(n19498), .op(n19500) );
  or2_1 U23528 ( .ip1(n24482), .ip2(n19498), .op(n19499) );
  nand2_1 U23529 ( .ip1(n19500), .ip2(n19499), .op(n19502) );
  nor2_1 U23530 ( .ip1(\x[49][6] ), .ip2(n23770), .op(n19501) );
  not_ab_or_c_or_d U23531 ( .ip1(sig_in[5]), .ip2(n19503), .ip3(n19502), .ip4(
        n19501), .op(n19505) );
  and2_1 U23532 ( .ip1(n24355), .ip2(\x[49][6] ), .op(n19504) );
  not_ab_or_c_or_d U23533 ( .ip1(\x[49][7] ), .ip2(n24044), .ip3(n19505), 
        .ip4(n19504), .op(n19506) );
  nor2_1 U23534 ( .ip1(n19507), .ip2(n19506), .op(n19632) );
  inv_1 U23535 ( .ip(n19632), .op(n19509) );
  nand2_1 U23536 ( .ip1(\x[49][8] ), .ip2(n23804), .op(n19508) );
  nand2_1 U23537 ( .ip1(n19509), .ip2(n19508), .op(n19512) );
  nor2_1 U23538 ( .ip1(\x[49][9] ), .ip2(n23981), .op(n19625) );
  or2_1 U23539 ( .ip1(n23779), .ip2(n19625), .op(n19511) );
  inv_1 U23540 ( .ip(\x[49][8] ), .op(n19626) );
  or2_1 U23541 ( .ip1(n19626), .ip2(n19625), .op(n19510) );
  nand2_1 U23542 ( .ip1(n19511), .ip2(n19510), .op(n19631) );
  nand2_1 U23543 ( .ip1(n19512), .ip2(n19631), .op(n19515) );
  and2_1 U23544 ( .ip1(n23146), .ip2(\x[49][10] ), .op(n19514) );
  not_ab_or_c_or_d U23545 ( .ip1(\x[49][9] ), .ip2(n24164), .ip3(n19514), 
        .ip4(n19513), .op(n19628) );
  nand2_1 U23546 ( .ip1(n19515), .ip2(n19628), .op(n19516) );
  nand2_1 U23547 ( .ip1(n19630), .ip2(n19516), .op(n19520) );
  inv_1 U23548 ( .ip(n19575), .op(n19517) );
  or2_1 U23549 ( .ip1(\x[49][12] ), .ip2(n19517), .op(n19519) );
  or2_1 U23550 ( .ip1(n24233), .ip2(n19517), .op(n19518) );
  nand2_1 U23551 ( .ip1(n19519), .ip2(n19518), .op(n19576) );
  nand2_1 U23552 ( .ip1(n19520), .ip2(n19576), .op(n19572) );
  nand2_1 U23553 ( .ip1(\x[48][15] ), .ip2(n24180), .op(n19523) );
  and2_1 U23554 ( .ip1(n23895), .ip2(\x[48][13] ), .op(n19521) );
  nor2_1 U23555 ( .ip1(\x[48][15] ), .ip2(n23143), .op(n19969) );
  not_ab_or_c_or_d U23556 ( .ip1(\x[48][14] ), .ip2(n24382), .ip3(n19521), 
        .ip4(n19969), .op(n19973) );
  nand2_1 U23557 ( .ip1(\x[48][12] ), .ip2(n24079), .op(n19522) );
  nand2_1 U23558 ( .ip1(n19973), .ip2(n19522), .op(n19964) );
  nand2_1 U23559 ( .ip1(n19523), .ip2(n19964), .op(n19571) );
  inv_1 U23560 ( .ip(n19523), .op(n19524) );
  or2_1 U23561 ( .ip1(sig_in[14]), .ip2(n19524), .op(n19527) );
  inv_1 U23562 ( .ip(\x[48][14] ), .op(n19525) );
  or2_1 U23563 ( .ip1(n19525), .ip2(n19524), .op(n19526) );
  nand2_1 U23564 ( .ip1(n19527), .ip2(n19526), .op(n19968) );
  nor2_1 U23565 ( .ip1(\x[48][13] ), .ip2(n24332), .op(n19528) );
  or2_1 U23566 ( .ip1(sig_in[12]), .ip2(n19528), .op(n19531) );
  inv_1 U23567 ( .ip(\x[48][12] ), .op(n19529) );
  or2_1 U23568 ( .ip1(n19529), .ip2(n19528), .op(n19530) );
  nand2_1 U23569 ( .ip1(n19531), .ip2(n19530), .op(n19965) );
  nor2_1 U23570 ( .ip1(\x[48][10] ), .ip2(n20880), .op(n19532) );
  or2_1 U23571 ( .ip1(sig_in[11]), .ip2(n19532), .op(n19535) );
  inv_1 U23572 ( .ip(\x[48][11] ), .op(n19533) );
  or2_1 U23573 ( .ip1(n19533), .ip2(n19532), .op(n19534) );
  nand2_1 U23574 ( .ip1(n19535), .ip2(n19534), .op(n19567) );
  inv_1 U23575 ( .ip(\x[48][7] ), .op(n19557) );
  nor2_1 U23576 ( .ip1(sig_in[7]), .ip2(n19557), .op(n19554) );
  inv_1 U23577 ( .ip(\x[48][5] ), .op(n19552) );
  nor2_1 U23578 ( .ip1(n22833), .ip2(n19552), .op(n19549) );
  inv_1 U23579 ( .ip(\x[48][3] ), .op(n19547) );
  and2_1 U23580 ( .ip1(n23659), .ip2(\x[48][2] ), .op(n19544) );
  inv_1 U23581 ( .ip(\x[48][1] ), .op(n19537) );
  inv_1 U23582 ( .ip(\x[48][0] ), .op(n19536) );
  not_ab_or_c_or_d U23583 ( .ip1(n24464), .ip2(n19537), .ip3(n23195), .ip4(
        n19536), .op(n19538) );
  or2_1 U23584 ( .ip1(\x[48][1] ), .ip2(n19538), .op(n19540) );
  or2_1 U23585 ( .ip1(n21685), .ip2(n19538), .op(n19539) );
  nand2_1 U23586 ( .ip1(n19540), .ip2(n19539), .op(n19542) );
  nor2_1 U23587 ( .ip1(\x[48][2] ), .ip2(n24463), .op(n19541) );
  nor2_1 U23588 ( .ip1(n19542), .ip2(n19541), .op(n19543) );
  not_ab_or_c_or_d U23589 ( .ip1(\x[48][3] ), .ip2(n24476), .ip3(n19544), 
        .ip4(n19543), .op(n19546) );
  nor2_1 U23590 ( .ip1(\x[48][4] ), .ip2(n23860), .op(n19545) );
  not_ab_or_c_or_d U23591 ( .ip1(n23251), .ip2(n19547), .ip3(n19546), .ip4(
        n19545), .op(n19548) );
  not_ab_or_c_or_d U23592 ( .ip1(\x[48][4] ), .ip2(n23860), .ip3(n19549), 
        .ip4(n19548), .op(n19551) );
  nor2_1 U23593 ( .ip1(\x[48][6] ), .ip2(n23770), .op(n19550) );
  not_ab_or_c_or_d U23594 ( .ip1(sig_in[5]), .ip2(n19552), .ip3(n19551), .ip4(
        n19550), .op(n19553) );
  not_ab_or_c_or_d U23595 ( .ip1(\x[48][6] ), .ip2(n24045), .ip3(n19554), 
        .ip4(n19553), .op(n19556) );
  nor2_1 U23596 ( .ip1(\x[48][8] ), .ip2(n24358), .op(n19555) );
  not_ab_or_c_or_d U23597 ( .ip1(n17732), .ip2(n19557), .ip3(n19556), .ip4(
        n19555), .op(n19558) );
  or2_1 U23598 ( .ip1(\x[48][8] ), .ip2(n19558), .op(n19560) );
  inv_1 U23599 ( .ip(sig_in[8]), .op(n24100) );
  or2_1 U23600 ( .ip1(n24100), .ip2(n19558), .op(n19559) );
  nand2_1 U23601 ( .ip1(n19560), .ip2(n19559), .op(n19562) );
  nor2_1 U23602 ( .ip1(\x[48][9] ), .ip2(n24269), .op(n19561) );
  or2_1 U23603 ( .ip1(n19562), .ip2(n19561), .op(n19565) );
  nand2_1 U23604 ( .ip1(\x[48][10] ), .ip2(n23146), .op(n19564) );
  nand2_1 U23605 ( .ip1(\x[48][9] ), .ip2(n24455), .op(n19563) );
  nand3_1 U23606 ( .ip1(n19565), .ip2(n19564), .ip3(n19563), .op(n19566) );
  nand2_1 U23607 ( .ip1(n19567), .ip2(n19566), .op(n19569) );
  inv_1 U23608 ( .ip(n17981), .op(n21793) );
  nand2_1 U23609 ( .ip1(\x[48][11] ), .ip2(n21793), .op(n19568) );
  nand2_1 U23610 ( .ip1(n19569), .ip2(n19568), .op(n19963) );
  nand3_1 U23611 ( .ip1(n19968), .ip2(n19965), .ip3(n19963), .op(n19570) );
  nand3_1 U23612 ( .ip1(n19572), .ip2(n19571), .ip3(n19570), .op(n19573) );
  not_ab_or_c_or_d U23613 ( .ip1(n19575), .ip2(n19636), .ip3(n19574), .ip4(
        n19573), .op(n24804) );
  inv_1 U23614 ( .ip(n19576), .op(n19641) );
  nor2_1 U23615 ( .ip1(\x[50][14] ), .ip2(n24230), .op(n19577) );
  or2_1 U23616 ( .ip1(\x[50][15] ), .ip2(n19577), .op(n19579) );
  or2_1 U23617 ( .ip1(n24384), .ip2(n19577), .op(n19578) );
  nand2_1 U23618 ( .ip1(n19579), .ip2(n19578), .op(n19624) );
  nand2_1 U23619 ( .ip1(\x[50][13] ), .ip2(n24235), .op(n19581) );
  nand2_1 U23620 ( .ip1(\x[50][14] ), .ip2(n24230), .op(n19580) );
  nand2_1 U23621 ( .ip1(n19581), .ip2(n19580), .op(n19623) );
  nor2_1 U23622 ( .ip1(\x[50][15] ), .ip2(n23143), .op(n19622) );
  not_ab_or_c_or_d U23623 ( .ip1(\x[50][11] ), .ip2(n24136), .ip3(\x[50][10] ), 
        .ip4(n24370), .op(n19614) );
  inv_1 U23624 ( .ip(\x[50][9] ), .op(n19606) );
  nor2_1 U23625 ( .ip1(\x[50][8] ), .ip2(n23971), .op(n19605) );
  and2_1 U23626 ( .ip1(n23804), .ip2(\x[50][8] ), .op(n19603) );
  inv_1 U23627 ( .ip(\x[50][6] ), .op(n19601) );
  nor2_1 U23628 ( .ip1(sig_in[6]), .ip2(n19601), .op(n19598) );
  nor2_1 U23629 ( .ip1(\x[50][3] ), .ip2(n24342), .op(n19591) );
  not_ab_or_c_or_d U23630 ( .ip1(\x[50][3] ), .ip2(n24476), .ip3(\x[50][2] ), 
        .ip4(n24470), .op(n19590) );
  nor2_1 U23631 ( .ip1(\x[50][4] ), .ip2(n24347), .op(n19589) );
  inv_1 U23632 ( .ip(\x[50][1] ), .op(n19583) );
  inv_1 U23633 ( .ip(\x[50][0] ), .op(n19582) );
  not_ab_or_c_or_d U23634 ( .ip1(n24464), .ip2(n19583), .ip3(sig_in[0]), .ip4(
        n19582), .op(n19587) );
  nand2_1 U23635 ( .ip1(\x[50][3] ), .ip2(n22525), .op(n19585) );
  nand2_1 U23636 ( .ip1(\x[50][1] ), .ip2(n21685), .op(n19584) );
  nand2_1 U23637 ( .ip1(n19585), .ip2(n19584), .op(n19586) );
  not_ab_or_c_or_d U23638 ( .ip1(\x[50][2] ), .ip2(n24107), .ip3(n19587), 
        .ip4(n19586), .op(n19588) );
  nor4_1 U23639 ( .ip1(n19591), .ip2(n19590), .ip3(n19589), .ip4(n19588), .op(
        n19592) );
  or2_1 U23640 ( .ip1(\x[50][4] ), .ip2(n19592), .op(n19594) );
  or2_1 U23641 ( .ip1(n23860), .ip2(n19592), .op(n19593) );
  nand2_1 U23642 ( .ip1(n19594), .ip2(n19593), .op(n19596) );
  nor2_1 U23643 ( .ip1(\x[50][5] ), .ip2(n24119), .op(n19595) );
  nor2_1 U23644 ( .ip1(n19596), .ip2(n19595), .op(n19597) );
  not_ab_or_c_or_d U23645 ( .ip1(\x[50][5] ), .ip2(n23600), .ip3(n19598), 
        .ip4(n19597), .op(n19600) );
  nor2_1 U23646 ( .ip1(\x[50][7] ), .ip2(n24142), .op(n19599) );
  not_ab_or_c_or_d U23647 ( .ip1(sig_in[6]), .ip2(n19601), .ip3(n19600), .ip4(
        n19599), .op(n19602) );
  not_ab_or_c_or_d U23648 ( .ip1(\x[50][7] ), .ip2(n24142), .ip3(n19603), 
        .ip4(n19602), .op(n19604) );
  not_ab_or_c_or_d U23649 ( .ip1(n21171), .ip2(n19606), .ip3(n19605), .ip4(
        n19604), .op(n19610) );
  nand2_1 U23650 ( .ip1(\x[50][11] ), .ip2(n21793), .op(n19608) );
  nand2_1 U23651 ( .ip1(\x[50][10] ), .ip2(n23146), .op(n19607) );
  nand2_1 U23652 ( .ip1(n19608), .ip2(n19607), .op(n19609) );
  not_ab_or_c_or_d U23653 ( .ip1(\x[50][9] ), .ip2(n24043), .ip3(n19610), 
        .ip4(n19609), .op(n19613) );
  nor2_1 U23654 ( .ip1(\x[50][11] ), .ip2(n21793), .op(n19612) );
  nor2_1 U23655 ( .ip1(\x[50][12] ), .ip2(n24079), .op(n19611) );
  or4_1 U23656 ( .ip1(n19614), .ip2(n19613), .ip3(n19612), .ip4(n19611), .op(
        n19616) );
  or2_1 U23657 ( .ip1(n24376), .ip2(\x[50][13] ), .op(n19615) );
  nand2_1 U23658 ( .ip1(n19624), .ip2(n19615), .op(n19617) );
  or2_1 U23659 ( .ip1(n19616), .ip2(n19617), .op(n19620) );
  nand2_1 U23660 ( .ip1(\x[50][12] ), .ip2(n24233), .op(n19618) );
  or2_1 U23661 ( .ip1(n19618), .ip2(n19617), .op(n19619) );
  nand2_1 U23662 ( .ip1(n19620), .ip2(n19619), .op(n19621) );
  not_ab_or_c_or_d U23663 ( .ip1(n19624), .ip2(n19623), .ip3(n19622), .ip4(
        n19621), .op(n19960) );
  or3_1 U23664 ( .ip1(sig_in[8]), .ip2(n19626), .ip3(n19625), .op(n19627) );
  nand2_1 U23665 ( .ip1(n19628), .ip2(n19627), .op(n19629) );
  nand2_1 U23666 ( .ip1(n19630), .ip2(n19629), .op(n19638) );
  nand3_1 U23667 ( .ip1(n19633), .ip2(n19632), .ip3(n19631), .op(n19637) );
  inv_1 U23668 ( .ip(n19634), .op(n19635) );
  not_ab_or_c_or_d U23669 ( .ip1(n19638), .ip2(n19637), .ip3(n19636), .ip4(
        n19635), .op(n19639) );
  not_ab_or_c_or_d U23670 ( .ip1(n19641), .ip2(n19640), .ip3(n19960), .ip4(
        n19639), .op(n24803) );
  nor2_1 U23671 ( .ip1(\x[52][14] ), .ip2(n24230), .op(n19642) );
  or2_1 U23672 ( .ip1(\x[52][15] ), .ip2(n19642), .op(n19644) );
  or2_1 U23673 ( .ip1(n24384), .ip2(n19642), .op(n19643) );
  nand2_1 U23674 ( .ip1(n19644), .ip2(n19643), .op(n19944) );
  nor2_1 U23675 ( .ip1(\x[52][15] ), .ip2(n23143), .op(n19686) );
  nor2_1 U23676 ( .ip1(n19944), .ip2(n19686), .op(n19945) );
  nor2_1 U23677 ( .ip1(\x[52][13] ), .ip2(n24081), .op(n19685) );
  nor2_1 U23678 ( .ip1(\x[52][12] ), .ip2(n24079), .op(n19684) );
  nor2_1 U23679 ( .ip1(\x[52][11] ), .ip2(n24456), .op(n19683) );
  and2_1 U23680 ( .ip1(n23146), .ip2(\x[52][10] ), .op(n19677) );
  inv_1 U23681 ( .ip(\x[52][9] ), .op(n19675) );
  nor2_1 U23682 ( .ip1(\x[52][8] ), .ip2(n24358), .op(n19674) );
  inv_1 U23683 ( .ip(\x[52][7] ), .op(n19667) );
  nor2_1 U23684 ( .ip1(sig_in[7]), .ip2(n19667), .op(n19665) );
  inv_1 U23685 ( .ip(\x[52][5] ), .op(n19663) );
  inv_1 U23686 ( .ip(\x[52][4] ), .op(n19655) );
  nor2_1 U23687 ( .ip1(n24462), .ip2(n19655), .op(n19653) );
  inv_1 U23688 ( .ip(\x[52][3] ), .op(n19651) );
  inv_1 U23689 ( .ip(\x[52][1] ), .op(n19646) );
  nor2_1 U23690 ( .ip1(n22513), .ip2(n19646), .op(n19648) );
  inv_1 U23691 ( .ip(\x[52][0] ), .op(n19645) );
  not_ab_or_c_or_d U23692 ( .ip1(n24464), .ip2(n19646), .ip3(n23195), .ip4(
        n19645), .op(n19647) );
  not_ab_or_c_or_d U23693 ( .ip1(\x[52][2] ), .ip2(n24107), .ip3(n19648), 
        .ip4(n19647), .op(n19650) );
  nor2_1 U23694 ( .ip1(\x[52][2] ), .ip2(n24463), .op(n19649) );
  not_ab_or_c_or_d U23695 ( .ip1(n24251), .ip2(n19651), .ip3(n19650), .ip4(
        n19649), .op(n19652) );
  not_ab_or_c_or_d U23696 ( .ip1(\x[52][3] ), .ip2(n22525), .ip3(n19653), 
        .ip4(n19652), .op(n19654) );
  or2_1 U23697 ( .ip1(sig_in[4]), .ip2(n19654), .op(n19657) );
  or2_1 U23698 ( .ip1(n19655), .ip2(n19654), .op(n19656) );
  nand2_1 U23699 ( .ip1(n19657), .ip2(n19656), .op(n19658) );
  or2_1 U23700 ( .ip1(\x[52][5] ), .ip2(n19658), .op(n19660) );
  or2_1 U23701 ( .ip1(n24482), .ip2(n19658), .op(n19659) );
  nand2_1 U23702 ( .ip1(n19660), .ip2(n19659), .op(n19662) );
  nor2_1 U23703 ( .ip1(\x[52][6] ), .ip2(n23770), .op(n19661) );
  not_ab_or_c_or_d U23704 ( .ip1(sig_in[5]), .ip2(n19663), .ip3(n19662), .ip4(
        n19661), .op(n19664) );
  not_ab_or_c_or_d U23705 ( .ip1(\x[52][6] ), .ip2(n24045), .ip3(n19665), 
        .ip4(n19664), .op(n19666) );
  or2_1 U23706 ( .ip1(n17732), .ip2(n19666), .op(n19669) );
  or2_1 U23707 ( .ip1(n19667), .ip2(n19666), .op(n19668) );
  nand2_1 U23708 ( .ip1(n19669), .ip2(n19668), .op(n19670) );
  or2_1 U23709 ( .ip1(\x[52][8] ), .ip2(n19670), .op(n19672) );
  or2_1 U23710 ( .ip1(n24100), .ip2(n19670), .op(n19671) );
  nand2_1 U23711 ( .ip1(n19672), .ip2(n19671), .op(n19673) );
  not_ab_or_c_or_d U23712 ( .ip1(n21171), .ip2(n19675), .ip3(n19674), .ip4(
        n19673), .op(n19676) );
  not_ab_or_c_or_d U23713 ( .ip1(\x[52][9] ), .ip2(n24164), .ip3(n19677), 
        .ip4(n19676), .op(n19679) );
  nor2_1 U23714 ( .ip1(n24370), .ip2(\x[52][10] ), .op(n19678) );
  nor2_1 U23715 ( .ip1(n19679), .ip2(n19678), .op(n19681) );
  and2_1 U23716 ( .ip1(n24371), .ip2(\x[52][11] ), .op(n19680) );
  nor2_1 U23717 ( .ip1(n19681), .ip2(n19680), .op(n19682) );
  nor4_1 U23718 ( .ip1(n19685), .ip2(n19684), .ip3(n19683), .ip4(n19682), .op(
        n19943) );
  inv_1 U23719 ( .ip(n19686), .op(n19690) );
  nand2_1 U23720 ( .ip1(\x[52][14] ), .ip2(n24327), .op(n19689) );
  nand2_1 U23721 ( .ip1(\x[52][12] ), .ip2(n24233), .op(n19688) );
  nand2_1 U23722 ( .ip1(\x[52][13] ), .ip2(n24081), .op(n19687) );
  nand4_1 U23723 ( .ip1(n19690), .ip2(n19689), .ip3(n19688), .ip4(n19687), 
        .op(n19946) );
  nor2_1 U23724 ( .ip1(n19943), .ip2(n19946), .op(n19733) );
  nor2_1 U23725 ( .ip1(n24239), .ip2(\x[51][11] ), .op(n19719) );
  and2_1 U23726 ( .ip1(n23146), .ip2(\x[51][10] ), .op(n19717) );
  inv_1 U23727 ( .ip(\x[51][9] ), .op(n19715) );
  and2_1 U23728 ( .ip1(n23804), .ip2(\x[51][8] ), .op(n19712) );
  inv_1 U23729 ( .ip(\x[51][7] ), .op(n19710) );
  nor2_1 U23730 ( .ip1(n17732), .ip2(n19710), .op(n19707) );
  inv_1 U23731 ( .ip(\x[51][3] ), .op(n19697) );
  inv_1 U23732 ( .ip(\x[51][1] ), .op(n19692) );
  nor2_1 U23733 ( .ip1(n22513), .ip2(n19692), .op(n19694) );
  inv_1 U23734 ( .ip(\x[51][0] ), .op(n19691) );
  not_ab_or_c_or_d U23735 ( .ip1(n24464), .ip2(n19692), .ip3(n23195), .ip4(
        n19691), .op(n19693) );
  not_ab_or_c_or_d U23736 ( .ip1(\x[51][2] ), .ip2(n24107), .ip3(n19694), 
        .ip4(n19693), .op(n19696) );
  nor2_1 U23737 ( .ip1(\x[51][2] ), .ip2(n23717), .op(n19695) );
  not_ab_or_c_or_d U23738 ( .ip1(n24251), .ip2(n19697), .ip3(n19696), .ip4(
        n19695), .op(n19701) );
  nand2_1 U23739 ( .ip1(\x[51][5] ), .ip2(n24119), .op(n19699) );
  nand2_1 U23740 ( .ip1(\x[51][4] ), .ip2(n23721), .op(n19698) );
  nand2_1 U23741 ( .ip1(n19699), .ip2(n19698), .op(n19700) );
  not_ab_or_c_or_d U23742 ( .ip1(\x[51][3] ), .ip2(n22525), .ip3(n19701), 
        .ip4(n19700), .op(n19705) );
  nor2_1 U23743 ( .ip1(\x[51][6] ), .ip2(n23770), .op(n19704) );
  nor2_1 U23744 ( .ip1(\x[51][5] ), .ip2(n24350), .op(n19703) );
  not_ab_or_c_or_d U23745 ( .ip1(\x[51][5] ), .ip2(n23600), .ip3(\x[51][4] ), 
        .ip4(n24347), .op(n19702) );
  nor4_1 U23746 ( .ip1(n19705), .ip2(n19704), .ip3(n19703), .ip4(n19702), .op(
        n19706) );
  not_ab_or_c_or_d U23747 ( .ip1(\x[51][6] ), .ip2(n24045), .ip3(n19707), 
        .ip4(n19706), .op(n19709) );
  nor2_1 U23748 ( .ip1(\x[51][8] ), .ip2(n24358), .op(n19708) );
  not_ab_or_c_or_d U23749 ( .ip1(n17732), .ip2(n19710), .ip3(n19709), .ip4(
        n19708), .op(n19711) );
  not_ab_or_c_or_d U23750 ( .ip1(\x[51][9] ), .ip2(n24043), .ip3(n19712), 
        .ip4(n19711), .op(n19714) );
  nor2_1 U23751 ( .ip1(\x[51][10] ), .ip2(n20880), .op(n19713) );
  not_ab_or_c_or_d U23752 ( .ip1(n21171), .ip2(n19715), .ip3(n19714), .ip4(
        n19713), .op(n19716) );
  not_ab_or_c_or_d U23753 ( .ip1(\x[51][11] ), .ip2(n24136), .ip3(n19717), 
        .ip4(n19716), .op(n19718) );
  or2_1 U23754 ( .ip1(n19719), .ip2(n19718), .op(n19953) );
  nor2_1 U23755 ( .ip1(\x[51][13] ), .ip2(n24376), .op(n19721) );
  nor2_1 U23756 ( .ip1(\x[51][12] ), .ip2(n24079), .op(n19720) );
  nor2_1 U23757 ( .ip1(n19721), .ip2(n19720), .op(n19955) );
  inv_1 U23758 ( .ip(n19955), .op(n19723) );
  nand2_1 U23759 ( .ip1(\x[51][15] ), .ip2(n24186), .op(n19728) );
  or2_1 U23760 ( .ip1(n24382), .ip2(\x[51][14] ), .op(n19722) );
  nand2_1 U23761 ( .ip1(n19728), .ip2(n19722), .op(n19952) );
  nor3_1 U23762 ( .ip1(n19953), .ip2(n19723), .ip3(n19952), .op(n19732) );
  nand2_1 U23763 ( .ip1(n24382), .ip2(\x[51][14] ), .op(n19725) );
  or2_1 U23764 ( .ip1(n24329), .ip2(\x[51][15] ), .op(n19951) );
  nand2_1 U23765 ( .ip1(\x[51][13] ), .ip2(n24081), .op(n19724) );
  nand3_1 U23766 ( .ip1(n19725), .ip2(n19951), .ip3(n19724), .op(n19957) );
  or2_1 U23767 ( .ip1(\x[51][12] ), .ip2(n19957), .op(n19727) );
  or2_1 U23768 ( .ip1(n24449), .ip2(n19957), .op(n19726) );
  nand2_1 U23769 ( .ip1(n19727), .ip2(n19726), .op(n19730) );
  inv_1 U23770 ( .ip(n19728), .op(n19729) );
  nor2_1 U23771 ( .ip1(n19730), .ip2(n19729), .op(n19731) );
  nor4_1 U23772 ( .ip1(n19945), .ip2(n19733), .ip3(n19732), .ip4(n19731), .op(
        n24821) );
  nor2_1 U23773 ( .ip1(\x[53][14] ), .ip2(n23938), .op(n19776) );
  inv_1 U23774 ( .ip(\x[53][12] ), .op(n19768) );
  nor2_1 U23775 ( .ip1(n19768), .ip2(n17845), .op(n19770) );
  inv_1 U23776 ( .ip(\x[53][8] ), .op(n19758) );
  and2_1 U23777 ( .ip1(n23659), .ip2(\x[53][2] ), .op(n19742) );
  inv_1 U23778 ( .ip(\x[53][1] ), .op(n19735) );
  inv_1 U23779 ( .ip(\x[53][0] ), .op(n19734) );
  not_ab_or_c_or_d U23780 ( .ip1(n24464), .ip2(n19735), .ip3(n23195), .ip4(
        n19734), .op(n19736) );
  or2_1 U23781 ( .ip1(\x[53][1] ), .ip2(n19736), .op(n19738) );
  or2_1 U23782 ( .ip1(n21685), .ip2(n19736), .op(n19737) );
  nand2_1 U23783 ( .ip1(n19738), .ip2(n19737), .op(n19740) );
  nor2_1 U23784 ( .ip1(\x[53][2] ), .ip2(n23717), .op(n19739) );
  nor2_1 U23785 ( .ip1(n19740), .ip2(n19739), .op(n19741) );
  not_ab_or_c_or_d U23786 ( .ip1(\x[53][3] ), .ip2(n22525), .ip3(n19742), 
        .ip4(n19741), .op(n19745) );
  nor2_1 U23787 ( .ip1(\x[53][5] ), .ip2(n24482), .op(n19746) );
  nor2_1 U23788 ( .ip1(\x[53][3] ), .ip2(n24342), .op(n19744) );
  nor2_1 U23789 ( .ip1(\x[53][4] ), .ip2(n23721), .op(n19743) );
  nor4_1 U23790 ( .ip1(n19745), .ip2(n19746), .ip3(n19744), .ip4(n19743), .op(
        n19752) );
  nand2_1 U23791 ( .ip1(n23600), .ip2(\x[53][5] ), .op(n19750) );
  inv_1 U23792 ( .ip(n19746), .op(n19747) );
  nand3_1 U23793 ( .ip1(\x[53][4] ), .ip2(n23721), .ip3(n19747), .op(n19749)
         );
  nand2_1 U23794 ( .ip1(\x[53][7] ), .ip2(n24044), .op(n19748) );
  nand3_1 U23795 ( .ip1(n19750), .ip2(n19749), .ip3(n19748), .op(n19751) );
  not_ab_or_c_or_d U23796 ( .ip1(\x[53][6] ), .ip2(n24045), .ip3(n19752), 
        .ip4(n19751), .op(n19756) );
  inv_1 U23797 ( .ip(\x[53][7] ), .op(n19754) );
  not_ab_or_c_or_d U23798 ( .ip1(\x[53][7] ), .ip2(n24492), .ip3(\x[53][6] ), 
        .ip4(n23770), .op(n19753) );
  nor2_1 U23799 ( .ip1(\x[53][9] ), .ip2(n23981), .op(n19757) );
  ab_or_c_or_d U23800 ( .ip1(n17732), .ip2(n19754), .ip3(n19753), .ip4(n19757), 
        .op(n19755) );
  not_ab_or_c_or_d U23801 ( .ip1(n23779), .ip2(n19758), .ip3(n19756), .ip4(
        n19755), .op(n19763) );
  nand2_1 U23802 ( .ip1(n20880), .ip2(\x[53][10] ), .op(n19761) );
  or3_1 U23803 ( .ip1(n19758), .ip2(n23779), .ip3(n19757), .op(n19760) );
  nand2_1 U23804 ( .ip1(\x[53][11] ), .ip2(n21793), .op(n19759) );
  nand3_1 U23805 ( .ip1(n19761), .ip2(n19760), .ip3(n19759), .op(n19762) );
  not_ab_or_c_or_d U23806 ( .ip1(\x[53][9] ), .ip2(n24164), .ip3(n19763), 
        .ip4(n19762), .op(n19767) );
  nor2_1 U23807 ( .ip1(n21793), .ip2(\x[53][11] ), .op(n19765) );
  not_ab_or_c_or_d U23808 ( .ip1(\x[53][11] ), .ip2(n24136), .ip3(\x[53][10] ), 
        .ip4(n20880), .op(n19764) );
  or2_1 U23809 ( .ip1(n19765), .ip2(n19764), .op(n19766) );
  not_ab_or_c_or_d U23810 ( .ip1(sig_in[12]), .ip2(n19768), .ip3(n19767), 
        .ip4(n19766), .op(n19769) );
  or2_1 U23811 ( .ip1(n19770), .ip2(n19769), .op(n19771) );
  or2_1 U23812 ( .ip1(\x[53][13] ), .ip2(n19771), .op(n19773) );
  or2_1 U23813 ( .ip1(n24137), .ip2(n19771), .op(n19772) );
  nand2_1 U23814 ( .ip1(n19773), .ip2(n19772), .op(n19775) );
  nor2_1 U23815 ( .ip1(\x[53][13] ), .ip2(n24137), .op(n19774) );
  nor3_1 U23816 ( .ip1(n19776), .ip2(n19775), .ip3(n19774), .op(n19780) );
  or2_1 U23817 ( .ip1(n24180), .ip2(\x[53][15] ), .op(n19778) );
  nand2_1 U23818 ( .ip1(\x[53][14] ), .ip2(n24327), .op(n19777) );
  nand2_1 U23819 ( .ip1(n19778), .ip2(n19777), .op(n19779) );
  nor2_1 U23820 ( .ip1(n19780), .ip2(n19779), .op(n19781) );
  or2_1 U23821 ( .ip1(\x[53][15] ), .ip2(n19781), .op(n19783) );
  or2_1 U23822 ( .ip1(n24329), .ip2(n19781), .op(n19782) );
  nand2_1 U23823 ( .ip1(n19783), .ip2(n19782), .op(n19949) );
  nor2_1 U23824 ( .ip1(\x[54][14] ), .ip2(n24230), .op(n19826) );
  nor2_1 U23825 ( .ip1(\x[54][11] ), .ip2(n24371), .op(n19820) );
  nor2_1 U23826 ( .ip1(\x[54][13] ), .ip2(n24081), .op(n19819) );
  nor2_1 U23827 ( .ip1(\x[54][12] ), .ip2(n24449), .op(n19818) );
  and2_1 U23828 ( .ip1(n23146), .ip2(\x[54][10] ), .op(n19812) );
  inv_1 U23829 ( .ip(\x[54][9] ), .op(n19810) );
  inv_1 U23830 ( .ip(\x[54][7] ), .op(n19802) );
  nor2_1 U23831 ( .ip1(n17732), .ip2(n19802), .op(n19800) );
  inv_1 U23832 ( .ip(\x[54][3] ), .op(n19790) );
  inv_1 U23833 ( .ip(\x[54][1] ), .op(n19785) );
  nor2_1 U23834 ( .ip1(n22513), .ip2(n19785), .op(n19787) );
  inv_1 U23835 ( .ip(\x[54][0] ), .op(n19784) );
  not_ab_or_c_or_d U23836 ( .ip1(sig_in[1]), .ip2(n19785), .ip3(sig_in[0]), 
        .ip4(n19784), .op(n19786) );
  not_ab_or_c_or_d U23837 ( .ip1(\x[54][2] ), .ip2(n24107), .ip3(n19787), 
        .ip4(n19786), .op(n19789) );
  nor2_1 U23838 ( .ip1(\x[54][2] ), .ip2(n23717), .op(n19788) );
  not_ab_or_c_or_d U23839 ( .ip1(n23251), .ip2(n19790), .ip3(n19789), .ip4(
        n19788), .op(n19794) );
  nand2_1 U23840 ( .ip1(\x[54][5] ), .ip2(n24119), .op(n19792) );
  nand2_1 U23841 ( .ip1(\x[54][4] ), .ip2(n23721), .op(n19791) );
  nand2_1 U23842 ( .ip1(n19792), .ip2(n19791), .op(n19793) );
  not_ab_or_c_or_d U23843 ( .ip1(\x[54][3] ), .ip2(n24476), .ip3(n19794), 
        .ip4(n19793), .op(n19798) );
  nor2_1 U23844 ( .ip1(\x[54][5] ), .ip2(n23283), .op(n19797) );
  nor2_1 U23845 ( .ip1(\x[54][6] ), .ip2(n23770), .op(n19796) );
  not_ab_or_c_or_d U23846 ( .ip1(\x[54][5] ), .ip2(n23600), .ip3(\x[54][4] ), 
        .ip4(n24347), .op(n19795) );
  nor4_1 U23847 ( .ip1(n19798), .ip2(n19797), .ip3(n19796), .ip4(n19795), .op(
        n19799) );
  not_ab_or_c_or_d U23848 ( .ip1(\x[54][6] ), .ip2(n24045), .ip3(n19800), 
        .ip4(n19799), .op(n19801) );
  or2_1 U23849 ( .ip1(n17732), .ip2(n19801), .op(n19804) );
  or2_1 U23850 ( .ip1(n19802), .ip2(n19801), .op(n19803) );
  nand2_1 U23851 ( .ip1(n19804), .ip2(n19803), .op(n19805) );
  or2_1 U23852 ( .ip1(\x[54][8] ), .ip2(n19805), .op(n19807) );
  or2_1 U23853 ( .ip1(n24491), .ip2(n19805), .op(n19806) );
  nand2_1 U23854 ( .ip1(n19807), .ip2(n19806), .op(n19809) );
  nor2_1 U23855 ( .ip1(\x[54][8] ), .ip2(n24358), .op(n19808) );
  not_ab_or_c_or_d U23856 ( .ip1(n21171), .ip2(n19810), .ip3(n19809), .ip4(
        n19808), .op(n19811) );
  not_ab_or_c_or_d U23857 ( .ip1(\x[54][9] ), .ip2(n24455), .ip3(n19812), 
        .ip4(n19811), .op(n19814) );
  nor2_1 U23858 ( .ip1(n23980), .ip2(\x[54][10] ), .op(n19813) );
  nor2_1 U23859 ( .ip1(n19814), .ip2(n19813), .op(n19816) );
  and2_1 U23860 ( .ip1(n24371), .ip2(\x[54][11] ), .op(n19815) );
  nor2_1 U23861 ( .ip1(n19816), .ip2(n19815), .op(n19817) );
  nor4_1 U23862 ( .ip1(n19820), .ip2(n19819), .ip3(n19818), .ip4(n19817), .op(
        n19824) );
  nand2_1 U23863 ( .ip1(\x[54][13] ), .ip2(n24081), .op(n19822) );
  nand2_1 U23864 ( .ip1(\x[54][12] ), .ip2(n24450), .op(n19821) );
  nand2_1 U23865 ( .ip1(n19822), .ip2(n19821), .op(n19823) );
  not_ab_or_c_or_d U23866 ( .ip1(\x[54][14] ), .ip2(n23938), .ip3(n19824), 
        .ip4(n19823), .op(n19825) );
  not_ab_or_c_or_d U23867 ( .ip1(\x[54][15] ), .ip2(n24384), .ip3(n19826), 
        .ip4(n19825), .op(n19827) );
  or2_1 U23868 ( .ip1(sig_in[15]), .ip2(n19827), .op(n19830) );
  inv_1 U23869 ( .ip(\x[54][15] ), .op(n19828) );
  or2_1 U23870 ( .ip1(n19828), .ip2(n19827), .op(n19829) );
  nand2_1 U23871 ( .ip1(n19830), .ip2(n19829), .op(n19875) );
  nor2_1 U23872 ( .ip1(n19949), .ip2(n19875), .op(n24824) );
  nor2_1 U23873 ( .ip1(\x[55][15] ), .ip2(n23143), .op(n19874) );
  nand2_1 U23874 ( .ip1(\x[55][13] ), .ip2(n24235), .op(n19832) );
  nand2_1 U23875 ( .ip1(\x[55][12] ), .ip2(n24079), .op(n19831) );
  nand2_1 U23876 ( .ip1(n19832), .ip2(n19831), .op(n19833) );
  not_ab_or_c_or_d U23877 ( .ip1(\x[55][14] ), .ip2(n24185), .ip3(n19874), 
        .ip4(n19833), .op(n19878) );
  inv_1 U23878 ( .ip(\x[55][12] ), .op(n19870) );
  nor2_1 U23879 ( .ip1(\x[55][13] ), .ip2(n24332), .op(n19869) );
  nor2_1 U23880 ( .ip1(\x[55][9] ), .ip2(n23981), .op(n19856) );
  inv_1 U23881 ( .ip(\x[55][8] ), .op(n19834) );
  nor3_1 U23882 ( .ip1(sig_in[8]), .ip2(n19856), .ip3(n19834), .op(n19860) );
  nor2_1 U23883 ( .ip1(\x[55][8] ), .ip2(n24358), .op(n19858) );
  nor2_1 U23884 ( .ip1(\x[55][7] ), .ip2(n24492), .op(n19857) );
  nor2_1 U23885 ( .ip1(\x[55][5] ), .ip2(n23600), .op(n19844) );
  inv_1 U23886 ( .ip(\x[55][4] ), .op(n19835) );
  nor3_1 U23887 ( .ip1(sig_in[4]), .ip2(n19844), .ip3(n19835), .op(n19847) );
  and2_1 U23888 ( .ip1(n23659), .ip2(\x[55][2] ), .op(n19841) );
  nand2_1 U23889 ( .ip1(\x[55][1] ), .ip2(n21685), .op(n19839) );
  nand2_1 U23890 ( .ip1(\x[55][0] ), .ip2(n24143), .op(n19838) );
  nor2_1 U23891 ( .ip1(\x[55][2] ), .ip2(n23717), .op(n19837) );
  nor2_1 U23892 ( .ip1(\x[55][1] ), .ip2(n21685), .op(n19836) );
  not_ab_or_c_or_d U23893 ( .ip1(n19839), .ip2(n19838), .ip3(n19837), .ip4(
        n19836), .op(n19840) );
  not_ab_or_c_or_d U23894 ( .ip1(\x[55][3] ), .ip2(n22525), .ip3(n19841), 
        .ip4(n19840), .op(n19845) );
  nor2_1 U23895 ( .ip1(\x[55][4] ), .ip2(n24256), .op(n19843) );
  nor2_1 U23896 ( .ip1(\x[55][3] ), .ip2(n24342), .op(n19842) );
  nor4_1 U23897 ( .ip1(n19845), .ip2(n19844), .ip3(n19843), .ip4(n19842), .op(
        n19846) );
  not_ab_or_c_or_d U23898 ( .ip1(\x[55][5] ), .ip2(n24482), .ip3(n19847), 
        .ip4(n19846), .op(n19849) );
  nor2_1 U23899 ( .ip1(\x[55][6] ), .ip2(n24355), .op(n19848) );
  or2_1 U23900 ( .ip1(n19849), .ip2(n19848), .op(n19851) );
  nand2_1 U23901 ( .ip1(\x[55][6] ), .ip2(n24485), .op(n19850) );
  nand2_1 U23902 ( .ip1(n19851), .ip2(n19850), .op(n19852) );
  or2_1 U23903 ( .ip1(\x[55][7] ), .ip2(n19852), .op(n19854) );
  or2_1 U23904 ( .ip1(n24142), .ip2(n19852), .op(n19853) );
  nand2_1 U23905 ( .ip1(n19854), .ip2(n19853), .op(n19855) );
  nor4_1 U23906 ( .ip1(n19858), .ip2(n19857), .ip3(n19856), .ip4(n19855), .op(
        n19859) );
  not_ab_or_c_or_d U23907 ( .ip1(\x[55][9] ), .ip2(n23981), .ip3(n19860), 
        .ip4(n19859), .op(n19864) );
  nand2_1 U23908 ( .ip1(\x[55][10] ), .ip2(n23146), .op(n19863) );
  nor2_1 U23909 ( .ip1(\x[55][10] ), .ip2(n20880), .op(n19862) );
  nor2_1 U23910 ( .ip1(\x[55][11] ), .ip2(n24239), .op(n19861) );
  not_ab_or_c_or_d U23911 ( .ip1(n19864), .ip2(n19863), .ip3(n19862), .ip4(
        n19861), .op(n19865) );
  or2_1 U23912 ( .ip1(\x[55][11] ), .ip2(n19865), .op(n19867) );
  or2_1 U23913 ( .ip1(n24239), .ip2(n19865), .op(n19866) );
  nand2_1 U23914 ( .ip1(n19867), .ip2(n19866), .op(n19868) );
  not_ab_or_c_or_d U23915 ( .ip1(sig_in[12]), .ip2(n19870), .ip3(n19869), 
        .ip4(n19868), .op(n19887) );
  inv_1 U23916 ( .ip(n19887), .op(n19877) );
  nor2_1 U23917 ( .ip1(\x[55][14] ), .ip2(n24185), .op(n19871) );
  or2_1 U23918 ( .ip1(\x[55][15] ), .ip2(n19871), .op(n19873) );
  or2_1 U23919 ( .ip1(n24384), .ip2(n19871), .op(n19872) );
  nand2_1 U23920 ( .ip1(n19873), .ip2(n19872), .op(n19886) );
  nor2_1 U23921 ( .ip1(n19886), .ip2(n19874), .op(n19879) );
  inv_1 U23922 ( .ip(n19875), .op(n19876) );
  not_ab_or_c_or_d U23923 ( .ip1(n19878), .ip2(n19877), .ip3(n19879), .ip4(
        n19876), .op(n24810) );
  nor2_1 U23924 ( .ip1(n19879), .ip2(n19878), .op(n19885) );
  nor2_1 U23925 ( .ip1(\x[56][15] ), .ip2(n23143), .op(n19928) );
  nand2_1 U23926 ( .ip1(n23143), .ip2(\x[56][15] ), .op(n19935) );
  inv_1 U23927 ( .ip(n19935), .op(n19880) );
  or2_1 U23928 ( .ip1(sig_in[14]), .ip2(n19880), .op(n19883) );
  inv_1 U23929 ( .ip(\x[56][14] ), .op(n19881) );
  or2_1 U23930 ( .ip1(n19881), .ip2(n19880), .op(n19882) );
  nand2_1 U23931 ( .ip1(n19883), .ip2(n19882), .op(n19937) );
  nor2_1 U23932 ( .ip1(n19928), .ip2(n19937), .op(n19884) );
  not_ab_or_c_or_d U23933 ( .ip1(n19887), .ip2(n19886), .ip3(n19885), .ip4(
        n19884), .op(n19932) );
  nand2_1 U23934 ( .ip1(\x[56][12] ), .ip2(n24233), .op(n19933) );
  nor2_1 U23935 ( .ip1(n24456), .ip2(\x[56][11] ), .op(n19889) );
  not_ab_or_c_or_d U23936 ( .ip1(\x[56][11] ), .ip2(n24239), .ip3(\x[56][10] ), 
        .ip4(n24370), .op(n19888) );
  or2_1 U23937 ( .ip1(n19889), .ip2(n19888), .op(n19921) );
  nor2_1 U23938 ( .ip1(\x[56][9] ), .ip2(n24455), .op(n19913) );
  nor2_1 U23939 ( .ip1(\x[56][7] ), .ip2(n24142), .op(n19912) );
  nor2_1 U23940 ( .ip1(\x[56][8] ), .ip2(n24491), .op(n19911) );
  nor2_1 U23941 ( .ip1(\x[56][5] ), .ip2(n24119), .op(n19899) );
  inv_1 U23942 ( .ip(\x[56][4] ), .op(n19890) );
  nor3_1 U23943 ( .ip1(n24462), .ip2(n19899), .ip3(n19890), .op(n19902) );
  and2_1 U23944 ( .ip1(n23659), .ip2(\x[56][2] ), .op(n19896) );
  inv_1 U23945 ( .ip(sig_in[1]), .op(n20652) );
  nand2_1 U23946 ( .ip1(\x[56][1] ), .ip2(n20652), .op(n19894) );
  nand2_1 U23947 ( .ip1(\x[56][0] ), .ip2(n24143), .op(n19893) );
  nor2_1 U23948 ( .ip1(\x[56][2] ), .ip2(n23717), .op(n19892) );
  nor2_1 U23949 ( .ip1(\x[56][1] ), .ip2(n20652), .op(n19891) );
  not_ab_or_c_or_d U23950 ( .ip1(n19894), .ip2(n19893), .ip3(n19892), .ip4(
        n19891), .op(n19895) );
  not_ab_or_c_or_d U23951 ( .ip1(\x[56][3] ), .ip2(n22525), .ip3(n19896), 
        .ip4(n19895), .op(n19900) );
  nor2_1 U23952 ( .ip1(\x[56][3] ), .ip2(n24342), .op(n19898) );
  nor2_1 U23953 ( .ip1(\x[56][4] ), .ip2(n24256), .op(n19897) );
  nor4_1 U23954 ( .ip1(n19900), .ip2(n19899), .ip3(n19898), .ip4(n19897), .op(
        n19901) );
  not_ab_or_c_or_d U23955 ( .ip1(\x[56][5] ), .ip2(n23600), .ip3(n19902), 
        .ip4(n19901), .op(n19904) );
  nor2_1 U23956 ( .ip1(\x[56][6] ), .ip2(n24485), .op(n19903) );
  or2_1 U23957 ( .ip1(n19904), .ip2(n19903), .op(n19906) );
  nand2_1 U23958 ( .ip1(\x[56][6] ), .ip2(n24485), .op(n19905) );
  nand2_1 U23959 ( .ip1(n19906), .ip2(n19905), .op(n19907) );
  or2_1 U23960 ( .ip1(\x[56][7] ), .ip2(n19907), .op(n19909) );
  or2_1 U23961 ( .ip1(n24142), .ip2(n19907), .op(n19908) );
  nand2_1 U23962 ( .ip1(n19909), .ip2(n19908), .op(n19910) );
  nor4_1 U23963 ( .ip1(n19913), .ip2(n19912), .ip3(n19911), .ip4(n19910), .op(
        n19919) );
  nand2_1 U23964 ( .ip1(\x[56][11] ), .ip2(n21793), .op(n19917) );
  inv_1 U23965 ( .ip(n19913), .op(n19914) );
  nand3_1 U23966 ( .ip1(\x[56][8] ), .ip2(n24491), .ip3(n19914), .op(n19916)
         );
  nand2_1 U23967 ( .ip1(\x[56][10] ), .ip2(n23146), .op(n19915) );
  nand3_1 U23968 ( .ip1(n19917), .ip2(n19916), .ip3(n19915), .op(n19918) );
  not_ab_or_c_or_d U23969 ( .ip1(\x[56][9] ), .ip2(n24043), .ip3(n19919), 
        .ip4(n19918), .op(n19920) );
  nor2_1 U23970 ( .ip1(n19921), .ip2(n19920), .op(n19939) );
  inv_1 U23971 ( .ip(n19939), .op(n19922) );
  nand2_1 U23972 ( .ip1(n19933), .ip2(n19922), .op(n19927) );
  buf_1 U23973 ( .ip(n24332), .op(n24137) );
  nor2_1 U23974 ( .ip1(\x[56][13] ), .ip2(n24137), .op(n19923) );
  or2_1 U23975 ( .ip1(sig_in[12]), .ip2(n19923), .op(n19926) );
  inv_1 U23976 ( .ip(\x[56][12] ), .op(n19924) );
  or2_1 U23977 ( .ip1(n19924), .ip2(n19923), .op(n19925) );
  nand2_1 U23978 ( .ip1(n19926), .ip2(n19925), .op(n19938) );
  nand2_1 U23979 ( .ip1(n19927), .ip2(n19938), .op(n19930) );
  and2_1 U23980 ( .ip1(n23895), .ip2(\x[56][13] ), .op(n19929) );
  not_ab_or_c_or_d U23981 ( .ip1(\x[56][14] ), .ip2(n24327), .ip3(n19929), 
        .ip4(n19928), .op(n19934) );
  nand2_1 U23982 ( .ip1(n19930), .ip2(n19934), .op(n19931) );
  nand2_1 U23983 ( .ip1(n19932), .ip2(n19931), .op(n24827) );
  nand2_1 U23984 ( .ip1(n19934), .ip2(n19933), .op(n19936) );
  nand2_1 U23985 ( .ip1(n19936), .ip2(n19935), .op(n19942) );
  nand3_1 U23986 ( .ip1(n19939), .ip2(n19938), .ip3(n19937), .op(n19940) );
  nand3_1 U23987 ( .ip1(n19942), .ip2(n19941), .ip3(n19940), .op(n24828) );
  nand2_1 U23988 ( .ip1(n24827), .ip2(n24828), .op(n24826) );
  nor3_1 U23989 ( .ip1(n24824), .ip2(n24810), .ip3(n24826), .op(n24807) );
  nand2_1 U23990 ( .ip1(n19944), .ip2(n19943), .op(n19950) );
  inv_1 U23991 ( .ip(n19945), .op(n19947) );
  nand2_1 U23992 ( .ip1(n19947), .ip2(n19946), .op(n19948) );
  nand3_1 U23993 ( .ip1(n19950), .ip2(n19949), .ip3(n19948), .op(n24809) );
  nand2_1 U23994 ( .ip1(n24807), .ip2(n24809), .op(n24822) );
  nor2_1 U23995 ( .ip1(n24821), .ip2(n24822), .op(n24840) );
  nand2_1 U23996 ( .ip1(n19952), .ip2(n19951), .op(n19962) );
  nand2_1 U23997 ( .ip1(\x[51][12] ), .ip2(n24449), .op(n19954) );
  nand2_1 U23998 ( .ip1(n19954), .ip2(n19953), .op(n19956) );
  nand2_1 U23999 ( .ip1(n19956), .ip2(n19955), .op(n19959) );
  inv_1 U24000 ( .ip(n19957), .op(n19958) );
  nand2_1 U24001 ( .ip1(n19959), .ip2(n19958), .op(n19961) );
  nand3_1 U24002 ( .ip1(n19962), .ip2(n19961), .ip3(n19960), .op(n24842) );
  nand2_1 U24003 ( .ip1(n24840), .ip2(n24842), .op(n24806) );
  nor3_1 U24004 ( .ip1(n24804), .ip2(n24803), .ip3(n24806), .op(n24816) );
  or2_1 U24005 ( .ip1(n19964), .ip2(n19963), .op(n19980) );
  inv_1 U24006 ( .ip(n19965), .op(n19972) );
  nor2_1 U24007 ( .ip1(n19967), .ip2(n19966), .op(n19971) );
  nor2_1 U24008 ( .ip1(n19969), .ip2(n19968), .op(n19970) );
  not_ab_or_c_or_d U24009 ( .ip1(n19973), .ip2(n19972), .ip3(n19971), .ip4(
        n19970), .op(n19979) );
  inv_1 U24010 ( .ip(n19974), .op(n19976) );
  nand3_1 U24011 ( .ip1(n19977), .ip2(n19976), .ip3(n19975), .op(n19978) );
  nand3_1 U24012 ( .ip1(n19980), .ip2(n19979), .ip3(n19978), .op(n24817) );
  nand2_1 U24013 ( .ip1(n24816), .ip2(n24817), .op(n24802) );
  nor2_1 U24014 ( .ip1(n24800), .ip2(n24802), .op(n24819) );
  nor2_1 U24015 ( .ip1(\x[45][15] ), .ip2(n23143), .op(n19984) );
  nor3_1 U24016 ( .ip1(n19984), .ip2(\x[45][14] ), .ip3(n24185), .op(n19981)
         );
  or2_1 U24017 ( .ip1(\x[45][15] ), .ip2(n19981), .op(n19983) );
  or2_1 U24018 ( .ip1(n24329), .ip2(n19981), .op(n19982) );
  nand2_1 U24019 ( .ip1(n19983), .ip2(n19982), .op(n20052) );
  nand2_1 U24020 ( .ip1(n24185), .ip2(\x[45][14] ), .op(n19987) );
  inv_1 U24021 ( .ip(n19984), .op(n19986) );
  nand2_1 U24022 ( .ip1(\x[45][13] ), .ip2(n24081), .op(n19985) );
  nand3_1 U24023 ( .ip1(n19987), .ip2(n19986), .ip3(n19985), .op(n20034) );
  or2_1 U24024 ( .ip1(\x[45][12] ), .ip2(n20034), .op(n19989) );
  or2_1 U24025 ( .ip1(n24233), .ip2(n20034), .op(n19988) );
  nand2_1 U24026 ( .ip1(n19989), .ip2(n19988), .op(n20047) );
  buf_1 U24027 ( .ip(n24137), .op(n24376) );
  or2_1 U24028 ( .ip1(\x[45][13] ), .ip2(n24376), .op(n19992) );
  inv_1 U24029 ( .ip(\x[45][12] ), .op(n19990) );
  nand2_1 U24030 ( .ip1(n17845), .ip2(n19990), .op(n19991) );
  nand2_1 U24031 ( .ip1(n19992), .ip2(n19991), .op(n20043) );
  inv_1 U24032 ( .ip(\x[45][11] ), .op(n20022) );
  nor2_1 U24033 ( .ip1(n20022), .ip2(n17981), .op(n20024) );
  and2_1 U24034 ( .ip1(n23146), .ip2(\x[45][10] ), .op(n20019) );
  inv_1 U24035 ( .ip(\x[45][9] ), .op(n20017) );
  nor2_1 U24036 ( .ip1(\x[45][8] ), .ip2(n24358), .op(n20016) );
  and2_1 U24037 ( .ip1(n24461), .ip2(\x[45][7] ), .op(n20009) );
  inv_1 U24038 ( .ip(\x[45][3] ), .op(n19999) );
  nor2_1 U24039 ( .ip1(\x[45][2] ), .ip2(n23717), .op(n19998) );
  inv_1 U24040 ( .ip(\x[45][1] ), .op(n19994) );
  nor2_1 U24041 ( .ip1(n22513), .ip2(n19994), .op(n19996) );
  inv_1 U24042 ( .ip(\x[45][0] ), .op(n19993) );
  not_ab_or_c_or_d U24043 ( .ip1(n24464), .ip2(n19994), .ip3(n23195), .ip4(
        n19993), .op(n19995) );
  not_ab_or_c_or_d U24044 ( .ip1(\x[45][2] ), .ip2(n24463), .ip3(n19996), 
        .ip4(n19995), .op(n19997) );
  not_ab_or_c_or_d U24045 ( .ip1(n23251), .ip2(n19999), .ip3(n19998), .ip4(
        n19997), .op(n20003) );
  nand2_1 U24046 ( .ip1(\x[45][5] ), .ip2(n24119), .op(n20001) );
  nand2_1 U24047 ( .ip1(\x[45][4] ), .ip2(n24256), .op(n20000) );
  nand2_1 U24048 ( .ip1(n20001), .ip2(n20000), .op(n20002) );
  not_ab_or_c_or_d U24049 ( .ip1(\x[45][3] ), .ip2(n24476), .ip3(n20003), 
        .ip4(n20002), .op(n20007) );
  nor2_1 U24050 ( .ip1(\x[45][6] ), .ip2(n24355), .op(n20006) );
  nor2_1 U24051 ( .ip1(\x[45][5] ), .ip2(n24350), .op(n20005) );
  not_ab_or_c_or_d U24052 ( .ip1(\x[45][5] ), .ip2(n24482), .ip3(\x[45][4] ), 
        .ip4(n24347), .op(n20004) );
  nor4_1 U24053 ( .ip1(n20007), .ip2(n20006), .ip3(n20005), .ip4(n20004), .op(
        n20008) );
  not_ab_or_c_or_d U24054 ( .ip1(\x[45][6] ), .ip2(n24045), .ip3(n20009), 
        .ip4(n20008), .op(n20011) );
  nor2_1 U24055 ( .ip1(\x[45][7] ), .ip2(n24142), .op(n20010) );
  nor2_1 U24056 ( .ip1(n20011), .ip2(n20010), .op(n20012) );
  or2_1 U24057 ( .ip1(\x[45][8] ), .ip2(n20012), .op(n20014) );
  or2_1 U24058 ( .ip1(n24100), .ip2(n20012), .op(n20013) );
  nand2_1 U24059 ( .ip1(n20014), .ip2(n20013), .op(n20015) );
  not_ab_or_c_or_d U24060 ( .ip1(sig_in[9]), .ip2(n20017), .ip3(n20016), .ip4(
        n20015), .op(n20018) );
  not_ab_or_c_or_d U24061 ( .ip1(\x[45][9] ), .ip2(n24164), .ip3(n20019), 
        .ip4(n20018), .op(n20021) );
  nor2_1 U24062 ( .ip1(\x[45][10] ), .ip2(n24457), .op(n20020) );
  not_ab_or_c_or_d U24063 ( .ip1(sig_in[11]), .ip2(n20022), .ip3(n20021), 
        .ip4(n20020), .op(n20023) );
  nor2_1 U24064 ( .ip1(n20024), .ip2(n20023), .op(n20048) );
  or2_1 U24065 ( .ip1(n20043), .ip2(n20048), .op(n20025) );
  nand2_1 U24066 ( .ip1(n20047), .ip2(n20025), .op(n20033) );
  and2_1 U24067 ( .ip1(n20027), .ip2(n20026), .op(n20032) );
  nor3_1 U24068 ( .ip1(n20030), .ip2(n20029), .ip3(n20028), .op(n20031) );
  ab_or_c_or_d U24069 ( .ip1(n20052), .ip2(n20033), .ip3(n20032), .ip4(n20031), 
        .op(n24838) );
  inv_1 U24070 ( .ip(n20034), .op(n20044) );
  inv_1 U24071 ( .ip(n20035), .op(n20038) );
  nor2_1 U24072 ( .ip1(n20036), .ip2(n20038), .op(n20042) );
  inv_1 U24073 ( .ip(n20037), .op(n20039) );
  nor3_1 U24074 ( .ip1(n20040), .ip2(n20039), .ip3(n20038), .op(n20041) );
  not_ab_or_c_or_d U24075 ( .ip1(n20044), .ip2(n20043), .ip3(n20042), .ip4(
        n20041), .op(n20051) );
  or2_1 U24076 ( .ip1(n20046), .ip2(n20045), .op(n20050) );
  nand2_1 U24077 ( .ip1(n20048), .ip2(n20047), .op(n20049) );
  nand4_1 U24078 ( .ip1(n20052), .ip2(n20051), .ip3(n20050), .ip4(n20049), 
        .op(n24820) );
  nand3_1 U24079 ( .ip1(n24819), .ip2(n24838), .ip3(n24820), .op(n24837) );
  nor2_1 U24080 ( .ip1(n24835), .ip2(n24837), .op(n25918) );
  nand2_1 U24081 ( .ip1(n26760), .ip2(n25918), .op(n27496) );
  nor3_1 U24082 ( .ip1(n24850), .ip2(n24852), .ip3(n27496), .op(n27533) );
  not_ab_or_c_or_d U24083 ( .ip1(n20056), .ip2(n20055), .ip3(n20054), .ip4(
        n20053), .op(n20058) );
  nor2_1 U24084 ( .ip1(n20058), .ip2(n20057), .op(n20110) );
  or2_1 U24085 ( .ip1(\x[71][14] ), .ip2(n20059), .op(n20061) );
  or2_1 U24086 ( .ip1(n23938), .ip2(n20059), .op(n20060) );
  nand2_1 U24087 ( .ip1(n20061), .ip2(n20060), .op(n20064) );
  inv_1 U24088 ( .ip(n20062), .op(n20063) );
  nor2_1 U24089 ( .ip1(n20064), .ip2(n20063), .op(n20109) );
  nand2_1 U24090 ( .ip1(n24384), .ip2(\x[72][15] ), .op(n20822) );
  inv_1 U24091 ( .ip(n20822), .op(n20065) );
  or2_1 U24092 ( .ip1(sig_in[14]), .ip2(n20065), .op(n20068) );
  inv_1 U24093 ( .ip(\x[72][14] ), .op(n20066) );
  or2_1 U24094 ( .ip1(n20066), .ip2(n20065), .op(n20067) );
  nand2_1 U24095 ( .ip1(n20068), .ip2(n20067), .op(n20836) );
  nor2_1 U24096 ( .ip1(\x[72][15] ), .ip2(n23143), .op(n20069) );
  nor2_1 U24097 ( .ip1(n20836), .ip2(n20069), .op(n20108) );
  and2_1 U24098 ( .ip1(n23895), .ip2(\x[72][13] ), .op(n20070) );
  not_ab_or_c_or_d U24099 ( .ip1(\x[72][14] ), .ip2(n24382), .ip3(n20070), 
        .ip4(n20069), .op(n20821) );
  nor2_1 U24100 ( .ip1(\x[72][13] ), .ip2(n24137), .op(n20072) );
  nor2_1 U24101 ( .ip1(\x[72][12] ), .ip2(n24449), .op(n20071) );
  nor2_1 U24102 ( .ip1(n20072), .ip2(n20071), .op(n20837) );
  inv_1 U24103 ( .ip(n20837), .op(n20073) );
  nand2_1 U24104 ( .ip1(n20821), .ip2(n20073), .op(n20106) );
  nand2_1 U24105 ( .ip1(\x[72][12] ), .ip2(n24450), .op(n20820) );
  inv_1 U24106 ( .ip(\x[72][11] ), .op(n20101) );
  and2_1 U24107 ( .ip1(n23146), .ip2(\x[72][10] ), .op(n20098) );
  inv_1 U24108 ( .ip(\x[72][9] ), .op(n20096) );
  and2_1 U24109 ( .ip1(n23804), .ip2(\x[72][8] ), .op(n20093) );
  nor2_1 U24110 ( .ip1(\x[72][5] ), .ip2(n24482), .op(n20083) );
  inv_1 U24111 ( .ip(\x[72][4] ), .op(n20074) );
  nor3_1 U24112 ( .ip1(n24462), .ip2(n20083), .ip3(n20074), .op(n20087) );
  nor2_1 U24113 ( .ip1(\x[72][4] ), .ip2(n23860), .op(n20085) );
  nor2_1 U24114 ( .ip1(\x[72][3] ), .ip2(n22525), .op(n20084) );
  nand2_1 U24115 ( .ip1(\x[72][1] ), .ip2(n20652), .op(n20077) );
  or2_1 U24116 ( .ip1(\x[72][1] ), .ip2(n20652), .op(n20075) );
  nand3_1 U24117 ( .ip1(n24143), .ip2(\x[72][0] ), .ip3(n20075), .op(n20076)
         );
  nand2_1 U24118 ( .ip1(n20077), .ip2(n20076), .op(n20079) );
  and2_1 U24119 ( .ip1(n22795), .ip2(\x[72][3] ), .op(n20078) );
  nor3_1 U24120 ( .ip1(\x[72][2] ), .ip2(n20079), .ip3(n20078), .op(n20081) );
  not_ab_or_c_or_d U24121 ( .ip1(n20079), .ip2(\x[72][2] ), .ip3(n20078), 
        .ip4(n24470), .op(n20080) );
  or2_1 U24122 ( .ip1(n20081), .ip2(n20080), .op(n20082) );
  nor4_1 U24123 ( .ip1(n20085), .ip2(n20084), .ip3(n20083), .ip4(n20082), .op(
        n20086) );
  not_ab_or_c_or_d U24124 ( .ip1(\x[72][5] ), .ip2(n23600), .ip3(n20087), 
        .ip4(n20086), .op(n20091) );
  nand2_1 U24125 ( .ip1(\x[72][6] ), .ip2(n24485), .op(n20090) );
  nor2_1 U24126 ( .ip1(\x[72][7] ), .ip2(n24044), .op(n20089) );
  nor2_1 U24127 ( .ip1(\x[72][6] ), .ip2(n24355), .op(n20088) );
  not_ab_or_c_or_d U24128 ( .ip1(n20091), .ip2(n20090), .ip3(n20089), .ip4(
        n20088), .op(n20092) );
  not_ab_or_c_or_d U24129 ( .ip1(\x[72][7] ), .ip2(n24044), .ip3(n20093), 
        .ip4(n20092), .op(n20095) );
  nor2_1 U24130 ( .ip1(\x[72][8] ), .ip2(n24491), .op(n20094) );
  not_ab_or_c_or_d U24131 ( .ip1(n21171), .ip2(n20096), .ip3(n20095), .ip4(
        n20094), .op(n20097) );
  not_ab_or_c_or_d U24132 ( .ip1(\x[72][9] ), .ip2(n24043), .ip3(n20098), 
        .ip4(n20097), .op(n20100) );
  nor2_1 U24133 ( .ip1(\x[72][10] ), .ip2(n20880), .op(n20099) );
  not_ab_or_c_or_d U24134 ( .ip1(sig_in[11]), .ip2(n20101), .ip3(n20100), 
        .ip4(n20099), .op(n20102) );
  or2_1 U24135 ( .ip1(\x[72][11] ), .ip2(n20102), .op(n20104) );
  or2_1 U24136 ( .ip1(n21793), .ip2(n20102), .op(n20103) );
  nand2_1 U24137 ( .ip1(n20104), .ip2(n20103), .op(n20834) );
  nand3_1 U24138 ( .ip1(n20821), .ip2(n20820), .ip3(n20834), .op(n20105) );
  nand2_1 U24139 ( .ip1(n20106), .ip2(n20105), .op(n20107) );
  nor4_1 U24140 ( .ip1(n20110), .ip2(n20109), .ip3(n20108), .ip4(n20107), .op(
        n24947) );
  nand2_1 U24141 ( .ip1(\x[74][15] ), .ip2(n24180), .op(n20201) );
  and2_1 U24142 ( .ip1(n23895), .ip2(\x[74][13] ), .op(n20111) );
  nor2_1 U24143 ( .ip1(\x[74][15] ), .ip2(n23143), .op(n20808) );
  not_ab_or_c_or_d U24144 ( .ip1(\x[74][14] ), .ip2(n24382), .ip3(n20111), 
        .ip4(n20808), .op(n20816) );
  nand2_1 U24145 ( .ip1(\x[74][12] ), .ip2(n24450), .op(n20813) );
  nand2_1 U24146 ( .ip1(n20816), .ip2(n20813), .op(n20200) );
  and2_1 U24147 ( .ip1(n24451), .ip2(\x[74][10] ), .op(n20114) );
  nor2_1 U24148 ( .ip1(\x[74][9] ), .ip2(n24164), .op(n20136) );
  inv_1 U24149 ( .ip(\x[74][8] ), .op(n20112) );
  nor3_1 U24150 ( .ip1(sig_in[8]), .ip2(n20136), .ip3(n20112), .op(n20113) );
  not_ab_or_c_or_d U24151 ( .ip1(\x[74][9] ), .ip2(n23981), .ip3(n20114), 
        .ip4(n20113), .op(n20117) );
  nor2_1 U24152 ( .ip1(\x[74][11] ), .ip2(n21793), .op(n20116) );
  nor2_1 U24153 ( .ip1(\x[74][10] ), .ip2(n20880), .op(n20115) );
  or2_1 U24154 ( .ip1(n20116), .ip2(n20115), .op(n20139) );
  or2_1 U24155 ( .ip1(n20117), .ip2(n20139), .op(n20142) );
  and2_1 U24156 ( .ip1(n24461), .ip2(\x[74][7] ), .op(n20134) );
  inv_1 U24157 ( .ip(\x[74][3] ), .op(n20124) );
  nor2_1 U24158 ( .ip1(\x[74][2] ), .ip2(n23717), .op(n20123) );
  inv_1 U24159 ( .ip(\x[74][1] ), .op(n20119) );
  nor2_1 U24160 ( .ip1(n22513), .ip2(n20119), .op(n20121) );
  inv_1 U24161 ( .ip(\x[74][0] ), .op(n20118) );
  not_ab_or_c_or_d U24162 ( .ip1(n24464), .ip2(n20119), .ip3(n23195), .ip4(
        n20118), .op(n20120) );
  not_ab_or_c_or_d U24163 ( .ip1(\x[74][2] ), .ip2(n24107), .ip3(n20121), 
        .ip4(n20120), .op(n20122) );
  not_ab_or_c_or_d U24164 ( .ip1(n23251), .ip2(n20124), .ip3(n20123), .ip4(
        n20122), .op(n20128) );
  nand2_1 U24165 ( .ip1(\x[74][5] ), .ip2(n24119), .op(n20126) );
  nand2_1 U24166 ( .ip1(\x[74][4] ), .ip2(n23721), .op(n20125) );
  nand2_1 U24167 ( .ip1(n20126), .ip2(n20125), .op(n20127) );
  not_ab_or_c_or_d U24168 ( .ip1(\x[74][3] ), .ip2(n24476), .ip3(n20128), 
        .ip4(n20127), .op(n20132) );
  nor2_1 U24169 ( .ip1(\x[74][5] ), .ip2(n23283), .op(n20131) );
  nor2_1 U24170 ( .ip1(\x[74][6] ), .ip2(n24355), .op(n20130) );
  not_ab_or_c_or_d U24171 ( .ip1(\x[74][5] ), .ip2(n24482), .ip3(\x[74][4] ), 
        .ip4(n24347), .op(n20129) );
  nor4_1 U24172 ( .ip1(n20132), .ip2(n20131), .ip3(n20130), .ip4(n20129), .op(
        n20133) );
  not_ab_or_c_or_d U24173 ( .ip1(\x[74][6] ), .ip2(n24045), .ip3(n20134), 
        .ip4(n20133), .op(n20138) );
  nor2_1 U24174 ( .ip1(\x[74][7] ), .ip2(n24044), .op(n20137) );
  nor2_1 U24175 ( .ip1(\x[74][8] ), .ip2(n24358), .op(n20135) );
  or4_1 U24176 ( .ip1(n20138), .ip2(n20137), .ip3(n20136), .ip4(n20135), .op(
        n20140) );
  or2_1 U24177 ( .ip1(n20140), .ip2(n20139), .op(n20141) );
  nand2_1 U24178 ( .ip1(n20142), .ip2(n20141), .op(n20143) );
  or2_1 U24179 ( .ip1(\x[74][11] ), .ip2(n20143), .op(n20145) );
  or2_1 U24180 ( .ip1(n24456), .ip2(n20143), .op(n20144) );
  nand2_1 U24181 ( .ip1(n20145), .ip2(n20144), .op(n20812) );
  nor2_1 U24182 ( .ip1(\x[74][13] ), .ip2(n24376), .op(n20147) );
  nor2_1 U24183 ( .ip1(\x[74][12] ), .ip2(n24449), .op(n20146) );
  nor2_1 U24184 ( .ip1(n20147), .ip2(n20146), .op(n20814) );
  inv_1 U24185 ( .ip(n20814), .op(n20149) );
  or2_1 U24186 ( .ip1(n24185), .ip2(\x[74][14] ), .op(n20148) );
  nand2_1 U24187 ( .ip1(n20201), .ip2(n20148), .op(n20807) );
  nor3_1 U24188 ( .ip1(n20812), .ip2(n20149), .ip3(n20807), .op(n20199) );
  and2_1 U24189 ( .ip1(n23895), .ip2(\x[75][13] ), .op(n20150) );
  nor2_1 U24190 ( .ip1(\x[75][15] ), .ip2(n23143), .op(n20156) );
  not_ab_or_c_or_d U24191 ( .ip1(\x[75][14] ), .ip2(n24185), .ip3(n20150), 
        .ip4(n20156), .op(n20197) );
  nor2_1 U24192 ( .ip1(\x[75][13] ), .ip2(n24137), .op(n20152) );
  nor2_1 U24193 ( .ip1(\x[75][12] ), .ip2(n24079), .op(n20151) );
  nor2_1 U24194 ( .ip1(n20152), .ip2(n20151), .op(n20756) );
  inv_1 U24195 ( .ip(n20756), .op(n20196) );
  nor2_1 U24196 ( .ip1(\x[75][14] ), .ip2(n23938), .op(n20153) );
  or2_1 U24197 ( .ip1(\x[75][15] ), .ip2(n20153), .op(n20155) );
  or2_1 U24198 ( .ip1(n24384), .ip2(n20153), .op(n20154) );
  nand2_1 U24199 ( .ip1(n20155), .ip2(n20154), .op(n20757) );
  nor2_1 U24200 ( .ip1(n20156), .ip2(n20757), .op(n20747) );
  inv_1 U24201 ( .ip(\x[75][7] ), .op(n20179) );
  nor2_1 U24202 ( .ip1(n17732), .ip2(n20179), .op(n20177) );
  inv_1 U24203 ( .ip(\x[75][5] ), .op(n20175) );
  inv_1 U24204 ( .ip(\x[75][4] ), .op(n20167) );
  nor2_1 U24205 ( .ip1(n24462), .ip2(n20167), .op(n20165) );
  inv_1 U24206 ( .ip(\x[75][3] ), .op(n20163) );
  inv_1 U24207 ( .ip(\x[75][1] ), .op(n20158) );
  nor2_1 U24208 ( .ip1(n22513), .ip2(n20158), .op(n20160) );
  inv_1 U24209 ( .ip(\x[75][0] ), .op(n20157) );
  not_ab_or_c_or_d U24210 ( .ip1(sig_in[1]), .ip2(n20158), .ip3(n23195), .ip4(
        n20157), .op(n20159) );
  not_ab_or_c_or_d U24211 ( .ip1(\x[75][2] ), .ip2(n24107), .ip3(n20160), 
        .ip4(n20159), .op(n20162) );
  nor2_1 U24212 ( .ip1(\x[75][2] ), .ip2(n23717), .op(n20161) );
  not_ab_or_c_or_d U24213 ( .ip1(n24251), .ip2(n20163), .ip3(n20162), .ip4(
        n20161), .op(n20164) );
  not_ab_or_c_or_d U24214 ( .ip1(\x[75][3] ), .ip2(n22525), .ip3(n20165), 
        .ip4(n20164), .op(n20166) );
  or2_1 U24215 ( .ip1(sig_in[4]), .ip2(n20166), .op(n20169) );
  or2_1 U24216 ( .ip1(n20167), .ip2(n20166), .op(n20168) );
  nand2_1 U24217 ( .ip1(n20169), .ip2(n20168), .op(n20170) );
  or2_1 U24218 ( .ip1(\x[75][5] ), .ip2(n20170), .op(n20172) );
  or2_1 U24219 ( .ip1(n23600), .ip2(n20170), .op(n20171) );
  nand2_1 U24220 ( .ip1(n20172), .ip2(n20171), .op(n20174) );
  nor2_1 U24221 ( .ip1(\x[75][6] ), .ip2(n24485), .op(n20173) );
  not_ab_or_c_or_d U24222 ( .ip1(sig_in[5]), .ip2(n20175), .ip3(n20174), .ip4(
        n20173), .op(n20176) );
  not_ab_or_c_or_d U24223 ( .ip1(\x[75][6] ), .ip2(n23509), .ip3(n20177), 
        .ip4(n20176), .op(n20178) );
  or2_1 U24224 ( .ip1(sig_in[7]), .ip2(n20178), .op(n20181) );
  or2_1 U24225 ( .ip1(n20179), .ip2(n20178), .op(n20180) );
  nand2_1 U24226 ( .ip1(n20181), .ip2(n20180), .op(n20182) );
  nand2_1 U24227 ( .ip1(\x[75][8] ), .ip2(n20182), .op(n20185) );
  nor2_1 U24228 ( .ip1(\x[75][9] ), .ip2(n24455), .op(n20184) );
  nor2_1 U24229 ( .ip1(\x[75][8] ), .ip2(n20182), .op(n20183) );
  ab_or_c_or_d U24230 ( .ip1(n23779), .ip2(n20185), .ip3(n20184), .ip4(n20183), 
        .op(n20189) );
  nand2_1 U24231 ( .ip1(\x[75][10] ), .ip2(n23146), .op(n20188) );
  nand2_1 U24232 ( .ip1(\x[75][11] ), .ip2(n21793), .op(n20187) );
  nand2_1 U24233 ( .ip1(\x[75][9] ), .ip2(n23981), .op(n20186) );
  and4_1 U24234 ( .ip1(n20189), .ip2(n20188), .ip3(n20187), .ip4(n20186), .op(
        n20193) );
  nor2_1 U24235 ( .ip1(n24371), .ip2(\x[75][11] ), .op(n20191) );
  not_ab_or_c_or_d U24236 ( .ip1(\x[75][11] ), .ip2(n24371), .ip3(\x[75][10] ), 
        .ip4(n20880), .op(n20190) );
  or2_1 U24237 ( .ip1(n20191), .ip2(n20190), .op(n20192) );
  nor2_1 U24238 ( .ip1(n20193), .ip2(n20192), .op(n20758) );
  nand2_1 U24239 ( .ip1(\x[75][12] ), .ip2(n24079), .op(n20194) );
  nand2_1 U24240 ( .ip1(n20197), .ip2(n20194), .op(n20746) );
  nor2_1 U24241 ( .ip1(n20758), .ip2(n20746), .op(n20195) );
  ab_or_c_or_d U24242 ( .ip1(n20197), .ip2(n20196), .ip3(n20747), .ip4(n20195), 
        .op(n20198) );
  not_ab_or_c_or_d U24243 ( .ip1(n20201), .ip2(n20200), .ip3(n20199), .ip4(
        n20198), .op(n24939) );
  and2_1 U24244 ( .ip1(n23895), .ip2(\x[76][13] ), .op(n20202) );
  nor2_1 U24245 ( .ip1(\x[76][15] ), .ip2(n23143), .op(n20751) );
  not_ab_or_c_or_d U24246 ( .ip1(\x[76][14] ), .ip2(n24230), .ip3(n20202), 
        .ip4(n20751), .op(n20755) );
  nand2_1 U24247 ( .ip1(\x[76][12] ), .ip2(n24450), .op(n20203) );
  nand2_1 U24248 ( .ip1(n20755), .ip2(n20203), .op(n20743) );
  nand2_1 U24249 ( .ip1(\x[76][15] ), .ip2(n24186), .op(n20293) );
  and2_1 U24250 ( .ip1(n23146), .ip2(\x[77][10] ), .op(n20204) );
  inv_1 U24251 ( .ip(\x[77][11] ), .op(n20206) );
  nor2_1 U24252 ( .ip1(n17981), .ip2(n20206), .op(n20209) );
  not_ab_or_c_or_d U24253 ( .ip1(\x[77][9] ), .ip2(n24269), .ip3(n20204), 
        .ip4(n20209), .op(n20718) );
  nor2_1 U24254 ( .ip1(\x[77][10] ), .ip2(n20880), .op(n20205) );
  or2_1 U24255 ( .ip1(sig_in[11]), .ip2(n20205), .op(n20208) );
  or2_1 U24256 ( .ip1(n20206), .ip2(n20205), .op(n20207) );
  nand2_1 U24257 ( .ip1(n20208), .ip2(n20207), .op(n20724) );
  nor2_1 U24258 ( .ip1(n20209), .ip2(n20724), .op(n20714) );
  or2_1 U24259 ( .ip1(n20718), .ip2(n20714), .op(n20239) );
  nor2_1 U24260 ( .ip1(\x[77][9] ), .ip2(n24455), .op(n20715) );
  or2_1 U24261 ( .ip1(n23779), .ip2(n20715), .op(n20211) );
  inv_1 U24262 ( .ip(\x[77][8] ), .op(n20716) );
  or2_1 U24263 ( .ip1(n20716), .ip2(n20715), .op(n20210) );
  nand2_1 U24264 ( .ip1(n20211), .ip2(n20210), .op(n20723) );
  nor2_1 U24265 ( .ip1(\x[77][5] ), .ip2(n23600), .op(n20224) );
  inv_1 U24266 ( .ip(\x[77][4] ), .op(n20212) );
  nor3_1 U24267 ( .ip1(sig_in[4]), .ip2(n20224), .ip3(n20212), .op(n20227) );
  and2_1 U24268 ( .ip1(n23659), .ip2(\x[77][2] ), .op(n20221) );
  inv_1 U24269 ( .ip(\x[77][1] ), .op(n20214) );
  inv_1 U24270 ( .ip(\x[77][0] ), .op(n20213) );
  not_ab_or_c_or_d U24271 ( .ip1(sig_in[1]), .ip2(n20214), .ip3(sig_in[0]), 
        .ip4(n20213), .op(n20215) );
  or2_1 U24272 ( .ip1(\x[77][1] ), .ip2(n20215), .op(n20217) );
  or2_1 U24273 ( .ip1(n20652), .ip2(n20215), .op(n20216) );
  nand2_1 U24274 ( .ip1(n20217), .ip2(n20216), .op(n20219) );
  nor2_1 U24275 ( .ip1(\x[77][2] ), .ip2(n23717), .op(n20218) );
  nor2_1 U24276 ( .ip1(n20219), .ip2(n20218), .op(n20220) );
  not_ab_or_c_or_d U24277 ( .ip1(\x[77][3] ), .ip2(n24476), .ip3(n20221), 
        .ip4(n20220), .op(n20225) );
  nor2_1 U24278 ( .ip1(\x[77][4] ), .ip2(n24347), .op(n20223) );
  nor2_1 U24279 ( .ip1(\x[77][3] ), .ip2(n24342), .op(n20222) );
  nor4_1 U24280 ( .ip1(n20225), .ip2(n20224), .ip3(n20223), .ip4(n20222), .op(
        n20226) );
  not_ab_or_c_or_d U24281 ( .ip1(\x[77][5] ), .ip2(n23600), .ip3(n20227), 
        .ip4(n20226), .op(n20231) );
  nand2_1 U24282 ( .ip1(\x[77][6] ), .ip2(n24045), .op(n20230) );
  nor2_1 U24283 ( .ip1(\x[77][6] ), .ip2(n23770), .op(n20229) );
  nor2_1 U24284 ( .ip1(\x[77][7] ), .ip2(n24142), .op(n20228) );
  not_ab_or_c_or_d U24285 ( .ip1(n20231), .ip2(n20230), .ip3(n20229), .ip4(
        n20228), .op(n20232) );
  or2_1 U24286 ( .ip1(\x[77][7] ), .ip2(n20232), .op(n20234) );
  or2_1 U24287 ( .ip1(n24461), .ip2(n20232), .op(n20233) );
  nand2_1 U24288 ( .ip1(n20234), .ip2(n20233), .op(n20721) );
  nand2_1 U24289 ( .ip1(\x[77][8] ), .ip2(n24100), .op(n20235) );
  nand2_1 U24290 ( .ip1(n20721), .ip2(n20235), .op(n20236) );
  nand2_1 U24291 ( .ip1(n20723), .ip2(n20236), .op(n20237) );
  or2_1 U24292 ( .ip1(n20237), .ip2(n20714), .op(n20238) );
  nand2_1 U24293 ( .ip1(n20239), .ip2(n20238), .op(n20242) );
  and2_1 U24294 ( .ip1(n23895), .ip2(\x[77][13] ), .op(n20240) );
  nor2_1 U24295 ( .ip1(\x[77][15] ), .ip2(n23143), .op(n20249) );
  not_ab_or_c_or_d U24296 ( .ip1(\x[77][14] ), .ip2(n23938), .ip3(n20240), 
        .ip4(n20249), .op(n20290) );
  nand2_1 U24297 ( .ip1(\x[77][12] ), .ip2(n24450), .op(n20241) );
  nand2_1 U24298 ( .ip1(n20290), .ip2(n20241), .op(n20733) );
  nor2_1 U24299 ( .ip1(n20242), .ip2(n20733), .op(n20292) );
  nor2_1 U24300 ( .ip1(\x[77][13] ), .ip2(n24376), .op(n20244) );
  nor2_1 U24301 ( .ip1(\x[77][12] ), .ip2(n24449), .op(n20243) );
  or2_1 U24302 ( .ip1(n20244), .ip2(n20243), .op(n20727) );
  nand2_1 U24303 ( .ip1(n23143), .ip2(\x[77][15] ), .op(n20732) );
  inv_1 U24304 ( .ip(n20732), .op(n20245) );
  or2_1 U24305 ( .ip1(sig_in[14]), .ip2(n20245), .op(n20248) );
  inv_1 U24306 ( .ip(\x[77][14] ), .op(n20246) );
  or2_1 U24307 ( .ip1(n20246), .ip2(n20245), .op(n20247) );
  nand2_1 U24308 ( .ip1(n20248), .ip2(n20247), .op(n20725) );
  nor2_1 U24309 ( .ip1(n20249), .ip2(n20725), .op(n20289) );
  inv_1 U24310 ( .ip(\x[76][11] ), .op(n20281) );
  and2_1 U24311 ( .ip1(n23146), .ip2(\x[76][10] ), .op(n20278) );
  inv_1 U24312 ( .ip(\x[76][9] ), .op(n20276) );
  nor2_1 U24313 ( .ip1(\x[76][8] ), .ip2(n24358), .op(n20275) );
  and2_1 U24314 ( .ip1(n24461), .ip2(\x[76][7] ), .op(n20268) );
  inv_1 U24315 ( .ip(\x[76][5] ), .op(n20266) );
  nor2_1 U24316 ( .ip1(n22833), .ip2(n20266), .op(n20263) );
  inv_1 U24317 ( .ip(\x[76][3] ), .op(n20261) );
  and2_1 U24318 ( .ip1(n24335), .ip2(\x[76][2] ), .op(n20258) );
  inv_1 U24319 ( .ip(\x[76][1] ), .op(n20251) );
  inv_1 U24320 ( .ip(\x[76][0] ), .op(n20250) );
  not_ab_or_c_or_d U24321 ( .ip1(sig_in[1]), .ip2(n20251), .ip3(n23195), .ip4(
        n20250), .op(n20252) );
  or2_1 U24322 ( .ip1(\x[76][1] ), .ip2(n20252), .op(n20254) );
  or2_1 U24323 ( .ip1(n21685), .ip2(n20252), .op(n20253) );
  nand2_1 U24324 ( .ip1(n20254), .ip2(n20253), .op(n20256) );
  nor2_1 U24325 ( .ip1(\x[76][2] ), .ip2(n23717), .op(n20255) );
  nor2_1 U24326 ( .ip1(n20256), .ip2(n20255), .op(n20257) );
  not_ab_or_c_or_d U24327 ( .ip1(\x[76][3] ), .ip2(n22525), .ip3(n20258), 
        .ip4(n20257), .op(n20260) );
  nor2_1 U24328 ( .ip1(\x[76][4] ), .ip2(n23721), .op(n20259) );
  not_ab_or_c_or_d U24329 ( .ip1(n24251), .ip2(n20261), .ip3(n20260), .ip4(
        n20259), .op(n20262) );
  not_ab_or_c_or_d U24330 ( .ip1(\x[76][4] ), .ip2(n23860), .ip3(n20263), 
        .ip4(n20262), .op(n20265) );
  nor2_1 U24331 ( .ip1(\x[76][6] ), .ip2(n23509), .op(n20264) );
  not_ab_or_c_or_d U24332 ( .ip1(sig_in[5]), .ip2(n20266), .ip3(n20265), .ip4(
        n20264), .op(n20267) );
  not_ab_or_c_or_d U24333 ( .ip1(\x[76][6] ), .ip2(n24045), .ip3(n20268), 
        .ip4(n20267), .op(n20270) );
  nor2_1 U24334 ( .ip1(\x[76][7] ), .ip2(n24492), .op(n20269) );
  nor2_1 U24335 ( .ip1(n20270), .ip2(n20269), .op(n20271) );
  or2_1 U24336 ( .ip1(\x[76][8] ), .ip2(n20271), .op(n20273) );
  or2_1 U24337 ( .ip1(n24100), .ip2(n20271), .op(n20272) );
  nand2_1 U24338 ( .ip1(n20273), .ip2(n20272), .op(n20274) );
  not_ab_or_c_or_d U24339 ( .ip1(n21171), .ip2(n20276), .ip3(n20275), .ip4(
        n20274), .op(n20277) );
  not_ab_or_c_or_d U24340 ( .ip1(\x[76][9] ), .ip2(n24043), .ip3(n20278), 
        .ip4(n20277), .op(n20280) );
  nor2_1 U24341 ( .ip1(\x[76][10] ), .ip2(n24457), .op(n20279) );
  not_ab_or_c_or_d U24342 ( .ip1(sig_in[11]), .ip2(n20281), .ip3(n20280), 
        .ip4(n20279), .op(n20282) );
  or2_1 U24343 ( .ip1(\x[76][11] ), .ip2(n20282), .op(n20284) );
  or2_1 U24344 ( .ip1(n24456), .ip2(n20282), .op(n20283) );
  nand2_1 U24345 ( .ip1(n20284), .ip2(n20283), .op(n20745) );
  nor2_1 U24346 ( .ip1(\x[76][13] ), .ip2(n24137), .op(n20286) );
  nor2_1 U24347 ( .ip1(\x[76][12] ), .ip2(n24079), .op(n20285) );
  or2_1 U24348 ( .ip1(n20286), .ip2(n20285), .op(n20754) );
  or2_1 U24349 ( .ip1(n24382), .ip2(\x[76][14] ), .op(n20287) );
  nand2_1 U24350 ( .ip1(n20293), .ip2(n20287), .op(n20749) );
  nor3_1 U24351 ( .ip1(n20745), .ip2(n20754), .ip3(n20749), .op(n20288) );
  ab_or_c_or_d U24352 ( .ip1(n20290), .ip2(n20727), .ip3(n20289), .ip4(n20288), 
        .op(n20291) );
  not_ab_or_c_or_d U24353 ( .ip1(n20743), .ip2(n20293), .ip3(n20292), .ip4(
        n20291), .op(n24648) );
  nor2_1 U24354 ( .ip1(\x[79][14] ), .ip2(n24230), .op(n20294) );
  or2_1 U24355 ( .ip1(\x[79][15] ), .ip2(n20294), .op(n20296) );
  or2_1 U24356 ( .ip1(n24329), .ip2(n20294), .op(n20295) );
  nand2_1 U24357 ( .ip1(n20296), .ip2(n20295), .op(n20704) );
  nor2_1 U24358 ( .ip1(\x[79][15] ), .ip2(n23143), .op(n20376) );
  nor2_1 U24359 ( .ip1(n20704), .ip2(n20376), .op(n20705) );
  nor2_1 U24360 ( .ip1(\x[78][13] ), .ip2(n24376), .op(n20297) );
  or2_1 U24361 ( .ip1(sig_in[12]), .ip2(n20297), .op(n20300) );
  inv_1 U24362 ( .ip(\x[78][12] ), .op(n20298) );
  or2_1 U24363 ( .ip1(n20298), .ip2(n20297), .op(n20299) );
  nand2_1 U24364 ( .ip1(n20300), .ip2(n20299), .op(n20737) );
  nor2_1 U24365 ( .ip1(\x[78][14] ), .ip2(n23938), .op(n20301) );
  or2_1 U24366 ( .ip1(\x[78][15] ), .ip2(n20301), .op(n20303) );
  or2_1 U24367 ( .ip1(n24329), .ip2(n20301), .op(n20302) );
  nand2_1 U24368 ( .ip1(n20303), .ip2(n20302), .op(n20336) );
  nor2_1 U24369 ( .ip1(\x[78][11] ), .ip2(n24456), .op(n20333) );
  and2_1 U24370 ( .ip1(n24451), .ip2(\x[78][10] ), .op(n20331) );
  nand2_1 U24371 ( .ip1(\x[78][7] ), .ip2(n24044), .op(n20324) );
  nand2_1 U24372 ( .ip1(\x[78][8] ), .ip2(n23971), .op(n20323) );
  nand2_1 U24373 ( .ip1(\x[78][9] ), .ip2(n23981), .op(n20322) );
  and2_1 U24374 ( .ip1(n23283), .ip2(\x[78][5] ), .op(n20312) );
  inv_1 U24375 ( .ip(\x[78][3] ), .op(n20310) );
  inv_1 U24376 ( .ip(\x[78][1] ), .op(n20305) );
  nor2_1 U24377 ( .ip1(n24464), .ip2(n20305), .op(n20307) );
  inv_1 U24378 ( .ip(\x[78][0] ), .op(n20304) );
  not_ab_or_c_or_d U24379 ( .ip1(sig_in[1]), .ip2(n20305), .ip3(n23195), .ip4(
        n20304), .op(n20306) );
  not_ab_or_c_or_d U24380 ( .ip1(\x[78][2] ), .ip2(n24107), .ip3(n20307), 
        .ip4(n20306), .op(n20309) );
  nor2_1 U24381 ( .ip1(\x[78][2] ), .ip2(n23717), .op(n20308) );
  not_ab_or_c_or_d U24382 ( .ip1(n24251), .ip2(n20310), .ip3(n20309), .ip4(
        n20308), .op(n20311) );
  not_ab_or_c_or_d U24383 ( .ip1(\x[78][3] ), .ip2(n22525), .ip3(n20312), 
        .ip4(n20311), .op(n20316) );
  nand2_1 U24384 ( .ip1(\x[78][4] ), .ip2(n23721), .op(n20315) );
  not_ab_or_c_or_d U24385 ( .ip1(\x[78][5] ), .ip2(n23600), .ip3(\x[78][4] ), 
        .ip4(n24347), .op(n20314) );
  nor2_1 U24386 ( .ip1(\x[78][5] ), .ip2(n24119), .op(n20313) );
  not_ab_or_c_or_d U24387 ( .ip1(n20316), .ip2(n20315), .ip3(n20314), .ip4(
        n20313), .op(n20317) );
  nand2_1 U24388 ( .ip1(n20317), .ip2(\x[78][6] ), .op(n20320) );
  nor2_1 U24389 ( .ip1(\x[78][7] ), .ip2(n24492), .op(n20319) );
  nor2_1 U24390 ( .ip1(n20317), .ip2(\x[78][6] ), .op(n20318) );
  ab_or_c_or_d U24391 ( .ip1(sig_in[6]), .ip2(n20320), .ip3(n20319), .ip4(
        n20318), .op(n20321) );
  and4_1 U24392 ( .ip1(n20324), .ip2(n20323), .ip3(n20322), .ip4(n20321), .op(
        n20328) );
  not_ab_or_c_or_d U24393 ( .ip1(\x[78][9] ), .ip2(n24043), .ip3(\x[78][8] ), 
        .ip4(n24358), .op(n20327) );
  nor2_1 U24394 ( .ip1(\x[78][10] ), .ip2(n20880), .op(n20326) );
  nor2_1 U24395 ( .ip1(\x[78][9] ), .ip2(n24455), .op(n20325) );
  nor4_1 U24396 ( .ip1(n20328), .ip2(n20327), .ip3(n20326), .ip4(n20325), .op(
        n20330) );
  and2_1 U24397 ( .ip1(n24371), .ip2(\x[78][11] ), .op(n20329) );
  nor3_1 U24398 ( .ip1(n20331), .ip2(n20330), .ip3(n20329), .op(n20332) );
  nor2_1 U24399 ( .ip1(n20333), .ip2(n20332), .op(n20734) );
  and3_1 U24400 ( .ip1(n20737), .ip2(n20336), .ip3(n20734), .op(n20383) );
  and2_1 U24401 ( .ip1(n23895), .ip2(\x[78][13] ), .op(n20334) );
  nor2_1 U24402 ( .ip1(\x[78][15] ), .ip2(n24090), .op(n20335) );
  not_ab_or_c_or_d U24403 ( .ip1(\x[78][14] ), .ip2(n24382), .ip3(n20334), 
        .ip4(n20335), .op(n20739) );
  nor2_1 U24404 ( .ip1(n20336), .ip2(n20335), .op(n20730) );
  or2_1 U24405 ( .ip1(n20739), .ip2(n20730), .op(n20338) );
  nand2_1 U24406 ( .ip1(\x[78][12] ), .ip2(n24450), .op(n20736) );
  or2_1 U24407 ( .ip1(n20736), .ip2(n20730), .op(n20337) );
  nand2_1 U24408 ( .ip1(n20338), .ip2(n20337), .op(n20382) );
  nor2_1 U24409 ( .ip1(\x[79][12] ), .ip2(n24079), .op(n20375) );
  nor2_1 U24410 ( .ip1(\x[79][11] ), .ip2(n24239), .op(n20374) );
  nor2_1 U24411 ( .ip1(\x[79][13] ), .ip2(n24137), .op(n20373) );
  and2_1 U24412 ( .ip1(n23146), .ip2(\x[79][10] ), .op(n20367) );
  inv_1 U24413 ( .ip(\x[79][9] ), .op(n20365) );
  and2_1 U24414 ( .ip1(n23804), .ip2(\x[79][8] ), .op(n20362) );
  inv_1 U24415 ( .ip(\x[79][6] ), .op(n20360) );
  nor2_1 U24416 ( .ip1(sig_in[6]), .ip2(n20360), .op(n20357) );
  inv_1 U24417 ( .ip(\x[79][3] ), .op(n20350) );
  and2_1 U24418 ( .ip1(n24335), .ip2(\x[79][2] ), .op(n20347) );
  inv_1 U24419 ( .ip(\x[79][1] ), .op(n20340) );
  inv_1 U24420 ( .ip(\x[79][0] ), .op(n20339) );
  not_ab_or_c_or_d U24421 ( .ip1(sig_in[1]), .ip2(n20340), .ip3(n23195), .ip4(
        n20339), .op(n20341) );
  or2_1 U24422 ( .ip1(\x[79][1] ), .ip2(n20341), .op(n20343) );
  or2_1 U24423 ( .ip1(n21685), .ip2(n20341), .op(n20342) );
  nand2_1 U24424 ( .ip1(n20343), .ip2(n20342), .op(n20345) );
  nor2_1 U24425 ( .ip1(\x[79][2] ), .ip2(n23717), .op(n20344) );
  nor2_1 U24426 ( .ip1(n20345), .ip2(n20344), .op(n20346) );
  not_ab_or_c_or_d U24427 ( .ip1(\x[79][3] ), .ip2(n24476), .ip3(n20347), 
        .ip4(n20346), .op(n20349) );
  nor2_1 U24428 ( .ip1(\x[79][4] ), .ip2(n24256), .op(n20348) );
  not_ab_or_c_or_d U24429 ( .ip1(n24251), .ip2(n20350), .ip3(n20349), .ip4(
        n20348), .op(n20351) );
  or2_1 U24430 ( .ip1(\x[79][4] ), .ip2(n20351), .op(n20353) );
  or2_1 U24431 ( .ip1(n23860), .ip2(n20351), .op(n20352) );
  nand2_1 U24432 ( .ip1(n20353), .ip2(n20352), .op(n20355) );
  nor2_1 U24433 ( .ip1(\x[79][5] ), .ip2(n24350), .op(n20354) );
  nor2_1 U24434 ( .ip1(n20355), .ip2(n20354), .op(n20356) );
  not_ab_or_c_or_d U24435 ( .ip1(\x[79][5] ), .ip2(n23600), .ip3(n20357), 
        .ip4(n20356), .op(n20359) );
  nor2_1 U24436 ( .ip1(\x[79][7] ), .ip2(n24492), .op(n20358) );
  not_ab_or_c_or_d U24437 ( .ip1(sig_in[6]), .ip2(n20360), .ip3(n20359), .ip4(
        n20358), .op(n20361) );
  not_ab_or_c_or_d U24438 ( .ip1(\x[79][7] ), .ip2(n24142), .ip3(n20362), 
        .ip4(n20361), .op(n20364) );
  nor2_1 U24439 ( .ip1(\x[79][8] ), .ip2(n24358), .op(n20363) );
  not_ab_or_c_or_d U24440 ( .ip1(sig_in[9]), .ip2(n20365), .ip3(n20364), .ip4(
        n20363), .op(n20366) );
  not_ab_or_c_or_d U24441 ( .ip1(\x[79][9] ), .ip2(n24455), .ip3(n20367), 
        .ip4(n20366), .op(n20369) );
  nor2_1 U24442 ( .ip1(n24370), .ip2(\x[79][10] ), .op(n20368) );
  nor2_1 U24443 ( .ip1(n20369), .ip2(n20368), .op(n20371) );
  and2_1 U24444 ( .ip1(n24239), .ip2(\x[79][11] ), .op(n20370) );
  nor2_1 U24445 ( .ip1(n20371), .ip2(n20370), .op(n20372) );
  nor4_1 U24446 ( .ip1(n20375), .ip2(n20374), .ip3(n20373), .ip4(n20372), .op(
        n20703) );
  nand2_1 U24447 ( .ip1(\x[79][12] ), .ip2(n24233), .op(n20380) );
  nand2_1 U24448 ( .ip1(\x[79][14] ), .ip2(n24327), .op(n20379) );
  nand2_1 U24449 ( .ip1(\x[79][13] ), .ip2(n24081), .op(n20378) );
  inv_1 U24450 ( .ip(n20376), .op(n20377) );
  nand4_1 U24451 ( .ip1(n20380), .ip2(n20379), .ip3(n20378), .ip4(n20377), 
        .op(n20707) );
  nor2_1 U24452 ( .ip1(n20703), .ip2(n20707), .op(n20381) );
  nor4_1 U24453 ( .ip1(n20705), .ip2(n20383), .ip3(n20382), .ip4(n20381), .op(
        n24925) );
  nor2_1 U24454 ( .ip1(\x[81][15] ), .ip2(n24090), .op(n20384) );
  or2_1 U24455 ( .ip1(\x[81][14] ), .ip2(n20384), .op(n20386) );
  or2_1 U24456 ( .ip1(n24382), .ip2(n20384), .op(n20385) );
  nand2_1 U24457 ( .ip1(n20386), .ip2(n20385), .op(n20469) );
  inv_1 U24458 ( .ip(\x[81][14] ), .op(n20389) );
  nor2_1 U24459 ( .ip1(\x[81][12] ), .ip2(n24079), .op(n20388) );
  nor2_1 U24460 ( .ip1(\x[81][13] ), .ip2(n24376), .op(n20387) );
  not_ab_or_c_or_d U24461 ( .ip1(sig_in[14]), .ip2(n20389), .ip3(n20388), 
        .ip4(n20387), .op(n20694) );
  inv_1 U24462 ( .ip(n20694), .op(n20468) );
  and2_1 U24463 ( .ip1(n24461), .ip2(\x[81][7] ), .op(n20403) );
  inv_1 U24464 ( .ip(\x[81][4] ), .op(n20401) );
  nor2_1 U24465 ( .ip1(n24462), .ip2(n20401), .op(n20398) );
  inv_1 U24466 ( .ip(\x[81][3] ), .op(n20396) );
  nor2_1 U24467 ( .ip1(\x[81][2] ), .ip2(n23717), .op(n20395) );
  inv_1 U24468 ( .ip(\x[81][1] ), .op(n20391) );
  nor2_1 U24469 ( .ip1(sig_in[1]), .ip2(n20391), .op(n20393) );
  inv_1 U24470 ( .ip(\x[81][0] ), .op(n20390) );
  not_ab_or_c_or_d U24471 ( .ip1(sig_in[1]), .ip2(n20391), .ip3(sig_in[0]), 
        .ip4(n20390), .op(n20392) );
  not_ab_or_c_or_d U24472 ( .ip1(\x[81][2] ), .ip2(n24107), .ip3(n20393), 
        .ip4(n20392), .op(n20394) );
  not_ab_or_c_or_d U24473 ( .ip1(n23251), .ip2(n20396), .ip3(n20395), .ip4(
        n20394), .op(n20397) );
  not_ab_or_c_or_d U24474 ( .ip1(\x[81][3] ), .ip2(n24476), .ip3(n20398), 
        .ip4(n20397), .op(n20400) );
  nor2_1 U24475 ( .ip1(\x[81][5] ), .ip2(n24482), .op(n20399) );
  not_ab_or_c_or_d U24476 ( .ip1(sig_in[4]), .ip2(n20401), .ip3(n20400), .ip4(
        n20399), .op(n20402) );
  not_ab_or_c_or_d U24477 ( .ip1(\x[81][5] ), .ip2(n24482), .ip3(n20403), 
        .ip4(n20402), .op(n20407) );
  nand2_1 U24478 ( .ip1(\x[81][6] ), .ip2(n24485), .op(n20406) );
  nor2_1 U24479 ( .ip1(\x[81][7] ), .ip2(n24142), .op(n20405) );
  not_ab_or_c_or_d U24480 ( .ip1(\x[81][7] ), .ip2(n24142), .ip3(\x[81][6] ), 
        .ip4(n23509), .op(n20404) );
  not_ab_or_c_or_d U24481 ( .ip1(n20407), .ip2(n20406), .ip3(n20405), .ip4(
        n20404), .op(n20408) );
  nand2_1 U24482 ( .ip1(\x[81][8] ), .ip2(n20408), .op(n20411) );
  nor2_1 U24483 ( .ip1(\x[81][9] ), .ip2(n24269), .op(n20410) );
  nor2_1 U24484 ( .ip1(\x[81][8] ), .ip2(n20408), .op(n20409) );
  ab_or_c_or_d U24485 ( .ip1(n23779), .ip2(n20411), .ip3(n20410), .ip4(n20409), 
        .op(n20415) );
  nand2_1 U24486 ( .ip1(\x[81][10] ), .ip2(n23146), .op(n20414) );
  nand2_1 U24487 ( .ip1(\x[81][11] ), .ip2(n21793), .op(n20413) );
  nand2_1 U24488 ( .ip1(\x[81][9] ), .ip2(n24043), .op(n20412) );
  and4_1 U24489 ( .ip1(n20415), .ip2(n20414), .ip3(n20413), .ip4(n20412), .op(
        n20419) );
  nor2_1 U24490 ( .ip1(n24239), .ip2(\x[81][11] ), .op(n20417) );
  not_ab_or_c_or_d U24491 ( .ip1(\x[81][11] ), .ip2(n24136), .ip3(\x[81][10] ), 
        .ip4(n24370), .op(n20416) );
  or2_1 U24492 ( .ip1(n20417), .ip2(n20416), .op(n20418) );
  nor2_1 U24493 ( .ip1(n20419), .ip2(n20418), .op(n20695) );
  nand2_1 U24494 ( .ip1(\x[81][12] ), .ip2(n24450), .op(n20421) );
  nand2_1 U24495 ( .ip1(\x[81][13] ), .ip2(n24235), .op(n20420) );
  nand3_1 U24496 ( .ip1(n20421), .ip2(n20469), .ip3(n20420), .op(n20696) );
  nor2_1 U24497 ( .ip1(n20695), .ip2(n20696), .op(n20467) );
  inv_1 U24498 ( .ip(\x[80][12] ), .op(n20463) );
  nor2_1 U24499 ( .ip1(\x[80][13] ), .ip2(n24137), .op(n20424) );
  or2_1 U24500 ( .ip1(n24382), .ip2(\x[80][14] ), .op(n20423) );
  nand2_1 U24501 ( .ip1(\x[80][15] ), .ip2(n24186), .op(n20422) );
  nand2_1 U24502 ( .ip1(n20423), .ip2(n20422), .op(n20464) );
  not_ab_or_c_or_d U24503 ( .ip1(sig_in[12]), .ip2(n20463), .ip3(n20424), 
        .ip4(n20464), .op(n20708) );
  nor2_1 U24504 ( .ip1(\x[80][15] ), .ip2(n24090), .op(n20459) );
  or2_1 U24505 ( .ip1(n20708), .ip2(n20459), .op(n20462) );
  inv_1 U24506 ( .ip(\x[80][9] ), .op(n20450) );
  not_ab_or_c_or_d U24507 ( .ip1(\x[80][9] ), .ip2(n24269), .ip3(\x[80][8] ), 
        .ip4(n24358), .op(n20449) );
  inv_1 U24508 ( .ip(\x[80][7] ), .op(n20443) );
  nor2_1 U24509 ( .ip1(n17732), .ip2(n20443), .op(n20441) );
  inv_1 U24510 ( .ip(\x[80][3] ), .op(n20431) );
  inv_1 U24511 ( .ip(\x[80][1] ), .op(n20426) );
  nor2_1 U24512 ( .ip1(n24464), .ip2(n20426), .op(n20428) );
  inv_1 U24513 ( .ip(\x[80][0] ), .op(n20425) );
  not_ab_or_c_or_d U24514 ( .ip1(sig_in[1]), .ip2(n20426), .ip3(n23195), .ip4(
        n20425), .op(n20427) );
  not_ab_or_c_or_d U24515 ( .ip1(\x[80][2] ), .ip2(n24335), .ip3(n20428), 
        .ip4(n20427), .op(n20430) );
  nor2_1 U24516 ( .ip1(\x[80][2] ), .ip2(n23717), .op(n20429) );
  not_ab_or_c_or_d U24517 ( .ip1(n24251), .ip2(n20431), .ip3(n20430), .ip4(
        n20429), .op(n20435) );
  nand2_1 U24518 ( .ip1(\x[80][5] ), .ip2(n23283), .op(n20433) );
  nand2_1 U24519 ( .ip1(\x[80][4] ), .ip2(n24347), .op(n20432) );
  nand2_1 U24520 ( .ip1(n20433), .ip2(n20432), .op(n20434) );
  not_ab_or_c_or_d U24521 ( .ip1(\x[80][3] ), .ip2(n22525), .ip3(n20435), 
        .ip4(n20434), .op(n20439) );
  nor2_1 U24522 ( .ip1(\x[80][5] ), .ip2(n23283), .op(n20438) );
  nor2_1 U24523 ( .ip1(\x[80][6] ), .ip2(n23509), .op(n20437) );
  not_ab_or_c_or_d U24524 ( .ip1(\x[80][5] ), .ip2(n23600), .ip3(\x[80][4] ), 
        .ip4(n24256), .op(n20436) );
  nor4_1 U24525 ( .ip1(n20439), .ip2(n20438), .ip3(n20437), .ip4(n20436), .op(
        n20440) );
  not_ab_or_c_or_d U24526 ( .ip1(\x[80][6] ), .ip2(n24045), .ip3(n20441), 
        .ip4(n20440), .op(n20442) );
  or2_1 U24527 ( .ip1(sig_in[7]), .ip2(n20442), .op(n20445) );
  or2_1 U24528 ( .ip1(n20443), .ip2(n20442), .op(n20444) );
  nand2_1 U24529 ( .ip1(n20445), .ip2(n20444), .op(n20447) );
  nor2_1 U24530 ( .ip1(n21171), .ip2(n20450), .op(n20446) );
  not_ab_or_c_or_d U24531 ( .ip1(\x[80][8] ), .ip2(n24100), .ip3(n20447), 
        .ip4(n20446), .op(n20448) );
  not_ab_or_c_or_d U24532 ( .ip1(sig_in[9]), .ip2(n20450), .ip3(n20449), .ip4(
        n20448), .op(n20451) );
  nand2_1 U24533 ( .ip1(\x[80][10] ), .ip2(n20451), .op(n20454) );
  nor2_1 U24534 ( .ip1(\x[80][11] ), .ip2(n24371), .op(n20453) );
  nor2_1 U24535 ( .ip1(\x[80][10] ), .ip2(n20451), .op(n20452) );
  ab_or_c_or_d U24536 ( .ip1(sig_in[10]), .ip2(n20454), .ip3(n20453), .ip4(
        n20452), .op(n20458) );
  nand2_1 U24537 ( .ip1(\x[80][14] ), .ip2(n23938), .op(n20457) );
  nand2_1 U24538 ( .ip1(\x[80][13] ), .ip2(n24235), .op(n20456) );
  nand2_1 U24539 ( .ip1(\x[80][11] ), .ip2(n21793), .op(n20455) );
  nand4_1 U24540 ( .ip1(n20458), .ip2(n20457), .ip3(n20456), .ip4(n20455), 
        .op(n20460) );
  or2_1 U24541 ( .ip1(n20460), .ip2(n20459), .op(n20461) );
  nand2_1 U24542 ( .ip1(n20462), .ip2(n20461), .op(n20710) );
  nand2_1 U24543 ( .ip1(\x[81][15] ), .ip2(n24186), .op(n20699) );
  or3_1 U24544 ( .ip1(n20464), .ip2(n20463), .ip3(n17845), .op(n20465) );
  nand3_1 U24545 ( .ip1(n20710), .ip2(n20699), .ip3(n20465), .op(n20466) );
  not_ab_or_c_or_d U24546 ( .ip1(n20469), .ip2(n20468), .ip3(n20467), .ip4(
        n20466), .op(n24910) );
  nor2_1 U24547 ( .ip1(\x[83][15] ), .ip2(n24090), .op(n20518) );
  nand2_1 U24548 ( .ip1(\x[83][13] ), .ip2(n24081), .op(n20471) );
  nand2_1 U24549 ( .ip1(\x[83][12] ), .ip2(n24449), .op(n20470) );
  nand2_1 U24550 ( .ip1(n20471), .ip2(n20470), .op(n20472) );
  not_ab_or_c_or_d U24551 ( .ip1(\x[83][14] ), .ip2(n24185), .ip3(n20518), 
        .ip4(n20472), .op(n20562) );
  nor2_1 U24552 ( .ip1(\x[83][10] ), .ip2(n24457), .op(n20473) );
  or2_1 U24553 ( .ip1(sig_in[11]), .ip2(n20473), .op(n20476) );
  inv_1 U24554 ( .ip(\x[83][11] ), .op(n20474) );
  or2_1 U24555 ( .ip1(n20474), .ip2(n20473), .op(n20475) );
  nand2_1 U24556 ( .ip1(n20476), .ip2(n20475), .op(n20510) );
  inv_1 U24557 ( .ip(\x[83][7] ), .op(n20500) );
  nor2_1 U24558 ( .ip1(sig_in[7]), .ip2(n20500), .op(n20497) );
  inv_1 U24559 ( .ip(\x[83][5] ), .op(n20495) );
  inv_1 U24560 ( .ip(\x[83][4] ), .op(n20487) );
  nor2_1 U24561 ( .ip1(n24462), .ip2(n20487), .op(n20485) );
  inv_1 U24562 ( .ip(\x[83][3] ), .op(n20483) );
  nor2_1 U24563 ( .ip1(\x[83][2] ), .ip2(n23717), .op(n20482) );
  inv_1 U24564 ( .ip(\x[83][1] ), .op(n20478) );
  nor2_1 U24565 ( .ip1(n24464), .ip2(n20478), .op(n20480) );
  inv_1 U24566 ( .ip(\x[83][0] ), .op(n20477) );
  not_ab_or_c_or_d U24567 ( .ip1(sig_in[1]), .ip2(n20478), .ip3(n23195), .ip4(
        n20477), .op(n20479) );
  not_ab_or_c_or_d U24568 ( .ip1(\x[83][2] ), .ip2(n23659), .ip3(n20480), 
        .ip4(n20479), .op(n20481) );
  not_ab_or_c_or_d U24569 ( .ip1(sig_in[3]), .ip2(n20483), .ip3(n20482), .ip4(
        n20481), .op(n20484) );
  not_ab_or_c_or_d U24570 ( .ip1(\x[83][3] ), .ip2(n24476), .ip3(n20485), 
        .ip4(n20484), .op(n20486) );
  or2_1 U24571 ( .ip1(sig_in[4]), .ip2(n20486), .op(n20489) );
  or2_1 U24572 ( .ip1(n20487), .ip2(n20486), .op(n20488) );
  nand2_1 U24573 ( .ip1(n20489), .ip2(n20488), .op(n20490) );
  or2_1 U24574 ( .ip1(\x[83][5] ), .ip2(n20490), .op(n20492) );
  or2_1 U24575 ( .ip1(n23600), .ip2(n20490), .op(n20491) );
  nand2_1 U24576 ( .ip1(n20492), .ip2(n20491), .op(n20494) );
  nor2_1 U24577 ( .ip1(\x[83][6] ), .ip2(n23509), .op(n20493) );
  not_ab_or_c_or_d U24578 ( .ip1(sig_in[5]), .ip2(n20495), .ip3(n20494), .ip4(
        n20493), .op(n20496) );
  not_ab_or_c_or_d U24579 ( .ip1(\x[83][6] ), .ip2(n24045), .ip3(n20497), 
        .ip4(n20496), .op(n20499) );
  nor2_1 U24580 ( .ip1(\x[83][8] ), .ip2(n24491), .op(n20498) );
  not_ab_or_c_or_d U24581 ( .ip1(n17732), .ip2(n20500), .ip3(n20499), .ip4(
        n20498), .op(n20501) );
  or2_1 U24582 ( .ip1(\x[83][8] ), .ip2(n20501), .op(n20503) );
  or2_1 U24583 ( .ip1(n24100), .ip2(n20501), .op(n20502) );
  nand2_1 U24584 ( .ip1(n20503), .ip2(n20502), .op(n20505) );
  nor2_1 U24585 ( .ip1(\x[83][9] ), .ip2(n24455), .op(n20504) );
  or2_1 U24586 ( .ip1(n20505), .ip2(n20504), .op(n20508) );
  nand2_1 U24587 ( .ip1(\x[83][10] ), .ip2(n23146), .op(n20507) );
  nand2_1 U24588 ( .ip1(\x[83][9] ), .ip2(n23981), .op(n20506) );
  nand3_1 U24589 ( .ip1(n20508), .ip2(n20507), .ip3(n20506), .op(n20509) );
  nand2_1 U24590 ( .ip1(n20510), .ip2(n20509), .op(n20514) );
  nand2_1 U24591 ( .ip1(\x[83][11] ), .ip2(n21793), .op(n20513) );
  nor2_1 U24592 ( .ip1(\x[83][12] ), .ip2(n24079), .op(n20512) );
  nor2_1 U24593 ( .ip1(\x[83][13] ), .ip2(n24376), .op(n20511) );
  not_ab_or_c_or_d U24594 ( .ip1(n20514), .ip2(n20513), .ip3(n20512), .ip4(
        n20511), .op(n20618) );
  inv_1 U24595 ( .ip(n20618), .op(n20561) );
  nor2_1 U24596 ( .ip1(\x[83][14] ), .ip2(n24230), .op(n20515) );
  or2_1 U24597 ( .ip1(\x[83][15] ), .ip2(n20515), .op(n20517) );
  or2_1 U24598 ( .ip1(n24180), .ip2(n20515), .op(n20516) );
  nand2_1 U24599 ( .ip1(n20517), .ip2(n20516), .op(n20619) );
  nor2_1 U24600 ( .ip1(n20619), .ip2(n20518), .op(n20563) );
  nor2_1 U24601 ( .ip1(n24384), .ip2(\x[82][15] ), .op(n20560) );
  and2_1 U24602 ( .ip1(n24332), .ip2(\x[82][13] ), .op(n20556) );
  inv_1 U24603 ( .ip(\x[82][12] ), .op(n20554) );
  nor2_1 U24604 ( .ip1(\x[82][11] ), .ip2(n24239), .op(n20548) );
  and2_1 U24605 ( .ip1(n24451), .ip2(\x[82][10] ), .op(n20546) );
  inv_1 U24606 ( .ip(\x[82][9] ), .op(n20543) );
  and2_1 U24607 ( .ip1(n23804), .ip2(\x[82][8] ), .op(n20540) );
  inv_1 U24608 ( .ip(\x[82][7] ), .op(n20538) );
  nor2_1 U24609 ( .ip1(n17732), .ip2(n20538), .op(n20535) );
  inv_1 U24610 ( .ip(\x[82][3] ), .op(n20525) );
  inv_1 U24611 ( .ip(\x[82][1] ), .op(n20520) );
  nor2_1 U24612 ( .ip1(n24464), .ip2(n20520), .op(n20522) );
  inv_1 U24613 ( .ip(\x[82][0] ), .op(n20519) );
  not_ab_or_c_or_d U24614 ( .ip1(sig_in[1]), .ip2(n20520), .ip3(n23195), .ip4(
        n20519), .op(n20521) );
  not_ab_or_c_or_d U24615 ( .ip1(\x[82][2] ), .ip2(n24107), .ip3(n20522), 
        .ip4(n20521), .op(n20524) );
  nor2_1 U24616 ( .ip1(\x[82][2] ), .ip2(n23717), .op(n20523) );
  not_ab_or_c_or_d U24617 ( .ip1(sig_in[3]), .ip2(n20525), .ip3(n20524), .ip4(
        n20523), .op(n20529) );
  nand2_1 U24618 ( .ip1(\x[82][5] ), .ip2(n24119), .op(n20527) );
  nand2_1 U24619 ( .ip1(\x[82][4] ), .ip2(n23721), .op(n20526) );
  nand2_1 U24620 ( .ip1(n20527), .ip2(n20526), .op(n20528) );
  not_ab_or_c_or_d U24621 ( .ip1(\x[82][3] ), .ip2(n22525), .ip3(n20529), 
        .ip4(n20528), .op(n20533) );
  nor2_1 U24622 ( .ip1(\x[82][6] ), .ip2(n23509), .op(n20532) );
  nor2_1 U24623 ( .ip1(\x[82][5] ), .ip2(n23600), .op(n20531) );
  not_ab_or_c_or_d U24624 ( .ip1(\x[82][5] ), .ip2(n24482), .ip3(\x[82][4] ), 
        .ip4(n24256), .op(n20530) );
  nor4_1 U24625 ( .ip1(n20533), .ip2(n20532), .ip3(n20531), .ip4(n20530), .op(
        n20534) );
  not_ab_or_c_or_d U24626 ( .ip1(\x[82][6] ), .ip2(n24045), .ip3(n20535), 
        .ip4(n20534), .op(n20537) );
  nor2_1 U24627 ( .ip1(\x[82][8] ), .ip2(n24491), .op(n20536) );
  not_ab_or_c_or_d U24628 ( .ip1(n17732), .ip2(n20538), .ip3(n20537), .ip4(
        n20536), .op(n20539) );
  not_ab_or_c_or_d U24629 ( .ip1(\x[82][9] ), .ip2(n24269), .ip3(n20540), 
        .ip4(n20539), .op(n20542) );
  nor2_1 U24630 ( .ip1(\x[82][10] ), .ip2(n24457), .op(n20541) );
  not_ab_or_c_or_d U24631 ( .ip1(sig_in[9]), .ip2(n20543), .ip3(n20542), .ip4(
        n20541), .op(n20545) );
  and2_1 U24632 ( .ip1(n24371), .ip2(\x[82][11] ), .op(n20544) );
  nor3_1 U24633 ( .ip1(n20546), .ip2(n20545), .ip3(n20544), .op(n20547) );
  nor2_1 U24634 ( .ip1(n20548), .ip2(n20547), .op(n20549) );
  or2_1 U24635 ( .ip1(\x[82][12] ), .ip2(n20549), .op(n20551) );
  or2_1 U24636 ( .ip1(n24449), .ip2(n20549), .op(n20550) );
  nand2_1 U24637 ( .ip1(n20551), .ip2(n20550), .op(n20553) );
  nor2_1 U24638 ( .ip1(\x[82][13] ), .ip2(n24137), .op(n20552) );
  not_ab_or_c_or_d U24639 ( .ip1(sig_in[12]), .ip2(n20554), .ip3(n20553), 
        .ip4(n20552), .op(n20555) );
  not_ab_or_c_or_d U24640 ( .ip1(\x[82][14] ), .ip2(n24382), .ip3(n20556), 
        .ip4(n20555), .op(n20558) );
  nor2_1 U24641 ( .ip1(\x[82][14] ), .ip2(n23938), .op(n20557) );
  not_ab_or_c_or_d U24642 ( .ip1(\x[82][15] ), .ip2(n24180), .ip3(n20558), 
        .ip4(n20557), .op(n20559) );
  or2_1 U24643 ( .ip1(n20560), .ip2(n20559), .op(n20702) );
  not_ab_or_c_or_d U24644 ( .ip1(n20562), .ip2(n20561), .ip3(n20563), .ip4(
        n20702), .op(n24913) );
  inv_1 U24645 ( .ip(n20562), .op(n20617) );
  inv_1 U24646 ( .ip(n20563), .op(n20616) );
  nor2_1 U24647 ( .ip1(\x[84][15] ), .ip2(n24090), .op(n20690) );
  and2_1 U24648 ( .ip1(n24186), .ip2(\x[84][15] ), .op(n20641) );
  or2_1 U24649 ( .ip1(sig_in[14]), .ip2(n20641), .op(n20566) );
  inv_1 U24650 ( .ip(\x[84][14] ), .op(n20564) );
  or2_1 U24651 ( .ip1(n20564), .ip2(n20641), .op(n20565) );
  nand2_1 U24652 ( .ip1(n20566), .ip2(n20565), .op(n20634) );
  nor2_1 U24653 ( .ip1(n20690), .ip2(n20634), .op(n20615) );
  nor2_1 U24654 ( .ip1(\x[84][13] ), .ip2(n24376), .op(n20567) );
  or2_1 U24655 ( .ip1(n17845), .ip2(n20567), .op(n20570) );
  inv_1 U24656 ( .ip(\x[84][12] ), .op(n20568) );
  or2_1 U24657 ( .ip1(n20568), .ip2(n20567), .op(n20569) );
  nand2_1 U24658 ( .ip1(n20570), .ip2(n20569), .op(n20633) );
  nand2_1 U24659 ( .ip1(n24079), .ip2(\x[84][12] ), .op(n20642) );
  inv_1 U24660 ( .ip(\x[84][11] ), .op(n20577) );
  nor2_1 U24661 ( .ip1(n20577), .ip2(n17981), .op(n20580) );
  and2_1 U24662 ( .ip1(\x[84][10] ), .ip2(n24451), .op(n20571) );
  nor2_1 U24663 ( .ip1(n20580), .ip2(n20571), .op(n20629) );
  inv_1 U24664 ( .ip(n20629), .op(n20572) );
  or2_1 U24665 ( .ip1(\x[84][9] ), .ip2(n20572), .op(n20574) );
  or2_1 U24666 ( .ip1(n24043), .ip2(n20572), .op(n20573) );
  nand2_1 U24667 ( .ip1(n20574), .ip2(n20573), .op(n20609) );
  nor2_1 U24668 ( .ip1(\x[84][9] ), .ip2(n24164), .op(n20628) );
  nor2_1 U24669 ( .ip1(\x[84][8] ), .ip2(n24491), .op(n20575) );
  nor2_1 U24670 ( .ip1(n20628), .ip2(n20575), .op(n20630) );
  inv_1 U24671 ( .ip(n20630), .op(n20608) );
  nor2_1 U24672 ( .ip1(\x[84][10] ), .ip2(n24457), .op(n20576) );
  or2_1 U24673 ( .ip1(sig_in[11]), .ip2(n20576), .op(n20579) );
  or2_1 U24674 ( .ip1(n20577), .ip2(n20576), .op(n20578) );
  nand2_1 U24675 ( .ip1(n20579), .ip2(n20578), .op(n20631) );
  nor2_1 U24676 ( .ip1(n20580), .ip2(n20631), .op(n20627) );
  inv_1 U24677 ( .ip(\x[84][7] ), .op(n20603) );
  nor2_1 U24678 ( .ip1(n17732), .ip2(n20603), .op(n20601) );
  inv_1 U24679 ( .ip(\x[84][5] ), .op(n20599) );
  nor2_1 U24680 ( .ip1(n22833), .ip2(n20599), .op(n20596) );
  inv_1 U24681 ( .ip(\x[84][3] ), .op(n20587) );
  inv_1 U24682 ( .ip(\x[84][1] ), .op(n20582) );
  nor2_1 U24683 ( .ip1(sig_in[1]), .ip2(n20582), .op(n20584) );
  inv_1 U24684 ( .ip(\x[84][0] ), .op(n20581) );
  not_ab_or_c_or_d U24685 ( .ip1(n24467), .ip2(n20582), .ip3(sig_in[0]), .ip4(
        n20581), .op(n20583) );
  not_ab_or_c_or_d U24686 ( .ip1(\x[84][2] ), .ip2(n24470), .ip3(n20584), 
        .ip4(n20583), .op(n20586) );
  nor2_1 U24687 ( .ip1(\x[84][2] ), .ip2(n23717), .op(n20585) );
  not_ab_or_c_or_d U24688 ( .ip1(sig_in[3]), .ip2(n20587), .ip3(n20586), .ip4(
        n20585), .op(n20588) );
  or2_1 U24689 ( .ip1(\x[84][3] ), .ip2(n20588), .op(n20590) );
  or2_1 U24690 ( .ip1(n22525), .ip2(n20588), .op(n20589) );
  nand2_1 U24691 ( .ip1(n20590), .ip2(n20589), .op(n20591) );
  or2_1 U24692 ( .ip1(sig_in[4]), .ip2(n20591), .op(n20594) );
  inv_1 U24693 ( .ip(\x[84][4] ), .op(n20592) );
  or2_1 U24694 ( .ip1(n20592), .ip2(n20591), .op(n20593) );
  nand2_1 U24695 ( .ip1(n20594), .ip2(n20593), .op(n20595) );
  not_ab_or_c_or_d U24696 ( .ip1(\x[84][4] ), .ip2(n24347), .ip3(n20596), 
        .ip4(n20595), .op(n20598) );
  nor2_1 U24697 ( .ip1(\x[84][6] ), .ip2(n23770), .op(n20597) );
  not_ab_or_c_or_d U24698 ( .ip1(n22833), .ip2(n20599), .ip3(n20598), .ip4(
        n20597), .op(n20600) );
  not_ab_or_c_or_d U24699 ( .ip1(\x[84][6] ), .ip2(n24045), .ip3(n20601), 
        .ip4(n20600), .op(n20602) );
  or2_1 U24700 ( .ip1(sig_in[7]), .ip2(n20602), .op(n20605) );
  or2_1 U24701 ( .ip1(n20603), .ip2(n20602), .op(n20604) );
  nand2_1 U24702 ( .ip1(n20605), .ip2(n20604), .op(n20632) );
  nand2_1 U24703 ( .ip1(\x[84][8] ), .ip2(n23971), .op(n20606) );
  nand2_1 U24704 ( .ip1(n20609), .ip2(n20606), .op(n20625) );
  nor2_1 U24705 ( .ip1(n20632), .ip2(n20625), .op(n20607) );
  ab_or_c_or_d U24706 ( .ip1(n20609), .ip2(n20608), .ip3(n20627), .ip4(n20607), 
        .op(n20610) );
  nand2_1 U24707 ( .ip1(n20642), .ip2(n20610), .op(n20613) );
  nand2_1 U24708 ( .ip1(\x[84][14] ), .ip2(n24327), .op(n20612) );
  nand2_1 U24709 ( .ip1(\x[84][13] ), .ip2(n24235), .op(n20611) );
  nand2_1 U24710 ( .ip1(n20612), .ip2(n20611), .op(n20639) );
  not_ab_or_c_or_d U24711 ( .ip1(n20633), .ip2(n20613), .ip3(n20690), .ip4(
        n20639), .op(n20614) );
  not_ab_or_c_or_d U24712 ( .ip1(n20617), .ip2(n20616), .ip3(n20615), .ip4(
        n20614), .op(n20621) );
  nand2_1 U24713 ( .ip1(n20619), .ip2(n20618), .op(n20620) );
  nand2_1 U24714 ( .ip1(n20621), .ip2(n20620), .op(n24919) );
  and2_1 U24715 ( .ip1(n24332), .ip2(\x[85][13] ), .op(n20622) );
  nor2_1 U24716 ( .ip1(\x[85][15] ), .ip2(n24180), .op(n20689) );
  not_ab_or_c_or_d U24717 ( .ip1(\x[85][14] ), .ip2(n24185), .ip3(n20622), 
        .ip4(n20689), .op(n20648) );
  nor2_1 U24718 ( .ip1(\x[85][13] ), .ip2(n24376), .op(n20624) );
  nor2_1 U24719 ( .ip1(\x[85][12] ), .ip2(n24449), .op(n20623) );
  nor2_1 U24720 ( .ip1(n20624), .ip2(n20623), .op(n20843) );
  inv_1 U24721 ( .ip(n20843), .op(n20647) );
  inv_1 U24722 ( .ip(n20625), .op(n20626) );
  ab_or_c_or_d U24723 ( .ip1(n20629), .ip2(n20628), .ip3(n20627), .ip4(n20626), 
        .op(n20638) );
  nand3_1 U24724 ( .ip1(n20632), .ip2(n20631), .ip3(n20630), .op(n20637) );
  inv_1 U24725 ( .ip(n20633), .op(n20636) );
  inv_1 U24726 ( .ip(n20634), .op(n20635) );
  not_ab_or_c_or_d U24727 ( .ip1(n20638), .ip2(n20637), .ip3(n20636), .ip4(
        n20635), .op(n20646) );
  inv_1 U24728 ( .ip(n20639), .op(n20640) );
  or2_1 U24729 ( .ip1(n20640), .ip2(n20641), .op(n20644) );
  or2_1 U24730 ( .ip1(n20642), .ip2(n20641), .op(n20643) );
  nand2_1 U24731 ( .ip1(n20644), .ip2(n20643), .op(n20645) );
  not_ab_or_c_or_d U24732 ( .ip1(n20648), .ip2(n20647), .ip3(n20646), .ip4(
        n20645), .op(n20693) );
  inv_1 U24733 ( .ip(n20648), .op(n20649) );
  or2_1 U24734 ( .ip1(\x[85][12] ), .ip2(n20649), .op(n20651) );
  or2_1 U24735 ( .ip1(n24079), .ip2(n20649), .op(n20650) );
  nand2_1 U24736 ( .ip1(n20651), .ip2(n20650), .op(n20841) );
  nor2_1 U24737 ( .ip1(n21793), .ip2(\x[85][11] ), .op(n20685) );
  inv_1 U24738 ( .ip(\x[85][5] ), .op(n20666) );
  nor2_1 U24739 ( .ip1(sig_in[5]), .ip2(n20666), .op(n20663) );
  inv_1 U24740 ( .ip(\x[85][3] ), .op(n20661) );
  and2_1 U24741 ( .ip1(n24335), .ip2(\x[85][2] ), .op(n20658) );
  nand2_1 U24742 ( .ip1(\x[85][1] ), .ip2(n20652), .op(n20656) );
  nand2_1 U24743 ( .ip1(\x[85][0] ), .ip2(n24143), .op(n20655) );
  nor2_1 U24744 ( .ip1(\x[85][2] ), .ip2(n23717), .op(n20654) );
  nor2_1 U24745 ( .ip1(\x[85][1] ), .ip2(n21685), .op(n20653) );
  not_ab_or_c_or_d U24746 ( .ip1(n20656), .ip2(n20655), .ip3(n20654), .ip4(
        n20653), .op(n20657) );
  not_ab_or_c_or_d U24747 ( .ip1(\x[85][3] ), .ip2(n22525), .ip3(n20658), 
        .ip4(n20657), .op(n20660) );
  nor2_1 U24748 ( .ip1(\x[85][4] ), .ip2(n23721), .op(n20659) );
  not_ab_or_c_or_d U24749 ( .ip1(sig_in[3]), .ip2(n20661), .ip3(n20660), .ip4(
        n20659), .op(n20662) );
  not_ab_or_c_or_d U24750 ( .ip1(\x[85][4] ), .ip2(n23860), .ip3(n20663), 
        .ip4(n20662), .op(n20665) );
  nor2_1 U24751 ( .ip1(\x[85][6] ), .ip2(n23770), .op(n20664) );
  not_ab_or_c_or_d U24752 ( .ip1(n22833), .ip2(n20666), .ip3(n20665), .ip4(
        n20664), .op(n20667) );
  or2_1 U24753 ( .ip1(\x[85][6] ), .ip2(n20667), .op(n20669) );
  or2_1 U24754 ( .ip1(n24045), .ip2(n20667), .op(n20668) );
  nand2_1 U24755 ( .ip1(n20669), .ip2(n20668), .op(n20670) );
  or2_1 U24756 ( .ip1(n17732), .ip2(n20670), .op(n20673) );
  inv_1 U24757 ( .ip(\x[85][7] ), .op(n20671) );
  or2_1 U24758 ( .ip1(n20671), .ip2(n20670), .op(n20672) );
  nand2_1 U24759 ( .ip1(n20673), .ip2(n20672), .op(n20677) );
  nand2_1 U24760 ( .ip1(\x[85][7] ), .ip2(n24492), .op(n20675) );
  nand2_1 U24761 ( .ip1(\x[85][9] ), .ip2(n24269), .op(n20674) );
  nand2_1 U24762 ( .ip1(n20675), .ip2(n20674), .op(n20676) );
  not_ab_or_c_or_d U24763 ( .ip1(\x[85][8] ), .ip2(n24100), .ip3(n20677), 
        .ip4(n20676), .op(n20681) );
  nor2_1 U24764 ( .ip1(\x[85][10] ), .ip2(n24457), .op(n20680) );
  not_ab_or_c_or_d U24765 ( .ip1(\x[85][9] ), .ip2(n24164), .ip3(\x[85][8] ), 
        .ip4(n24358), .op(n20679) );
  nor2_1 U24766 ( .ip1(\x[85][9] ), .ip2(n24455), .op(n20678) );
  nor4_1 U24767 ( .ip1(n20681), .ip2(n20680), .ip3(n20679), .ip4(n20678), .op(
        n20683) );
  and2_1 U24768 ( .ip1(n24451), .ip2(\x[85][10] ), .op(n20682) );
  not_ab_or_c_or_d U24769 ( .ip1(\x[85][11] ), .ip2(n24136), .ip3(n20683), 
        .ip4(n20682), .op(n20684) );
  nor2_1 U24770 ( .ip1(n20685), .ip2(n20684), .op(n20845) );
  inv_1 U24771 ( .ip(n20845), .op(n20691) );
  nor2_1 U24772 ( .ip1(\x[85][14] ), .ip2(n23938), .op(n20686) );
  or2_1 U24773 ( .ip1(\x[85][15] ), .ip2(n20686), .op(n20688) );
  or2_1 U24774 ( .ip1(n24384), .ip2(n20686), .op(n20687) );
  nand2_1 U24775 ( .ip1(n20688), .ip2(n20687), .op(n20844) );
  nor2_1 U24776 ( .ip1(n20689), .ip2(n20844), .op(n20842) );
  not_ab_or_c_or_d U24777 ( .ip1(n20841), .ip2(n20691), .ip3(n20690), .ip4(
        n20842), .op(n20692) );
  nand2_1 U24778 ( .ip1(n20693), .ip2(n20692), .op(n24920) );
  nand2_1 U24779 ( .ip1(n24919), .ip2(n24920), .op(n24915) );
  nor2_1 U24780 ( .ip1(n24913), .ip2(n24915), .op(n24916) );
  nand2_1 U24781 ( .ip1(n20695), .ip2(n20694), .op(n20698) );
  inv_1 U24782 ( .ip(n20696), .op(n20697) );
  nand2_1 U24783 ( .ip1(n20698), .ip2(n20697), .op(n20700) );
  nand2_1 U24784 ( .ip1(n20700), .ip2(n20699), .op(n20701) );
  nand2_1 U24785 ( .ip1(n20702), .ip2(n20701), .op(n24917) );
  nand2_1 U24786 ( .ip1(n24916), .ip2(n24917), .op(n24912) );
  nor2_1 U24787 ( .ip1(n24910), .ip2(n24912), .op(n24928) );
  nand2_1 U24788 ( .ip1(n20704), .ip2(n20703), .op(n20713) );
  inv_1 U24789 ( .ip(n20705), .op(n20706) );
  nand2_1 U24790 ( .ip1(n20707), .ip2(n20706), .op(n20712) );
  nand3_1 U24791 ( .ip1(n24233), .ip2(n20708), .ip3(\x[80][12] ), .op(n20709)
         );
  nand2_1 U24792 ( .ip1(n20710), .ip2(n20709), .op(n20711) );
  nand3_1 U24793 ( .ip1(n20713), .ip2(n20712), .ip3(n20711), .op(n24929) );
  nand2_1 U24794 ( .ip1(n24928), .ip2(n24929), .op(n24927) );
  nor2_1 U24795 ( .ip1(n24925), .ip2(n24927), .op(n24931) );
  inv_1 U24796 ( .ip(n20714), .op(n20720) );
  or3_1 U24797 ( .ip1(sig_in[8]), .ip2(n20716), .ip3(n20715), .op(n20717) );
  nand2_1 U24798 ( .ip1(n20718), .ip2(n20717), .op(n20719) );
  nand2_1 U24799 ( .ip1(n20720), .ip2(n20719), .op(n20729) );
  inv_1 U24800 ( .ip(n20721), .op(n20722) );
  nand3_1 U24801 ( .ip1(n20724), .ip2(n20723), .ip3(n20722), .op(n20728) );
  inv_1 U24802 ( .ip(n20725), .op(n20726) );
  not_ab_or_c_or_d U24803 ( .ip1(n20729), .ip2(n20728), .ip3(n20727), .ip4(
        n20726), .op(n20731) );
  not_ab_or_c_or_d U24804 ( .ip1(n20733), .ip2(n20732), .ip3(n20731), .ip4(
        n20730), .op(n20742) );
  inv_1 U24805 ( .ip(n20734), .op(n20735) );
  nand2_1 U24806 ( .ip1(n20736), .ip2(n20735), .op(n20738) );
  nand2_1 U24807 ( .ip1(n20738), .ip2(n20737), .op(n20740) );
  nand2_1 U24808 ( .ip1(n20740), .ip2(n20739), .op(n20741) );
  nand2_1 U24809 ( .ip1(n20742), .ip2(n20741), .op(n24933) );
  nand2_1 U24810 ( .ip1(n24931), .ip2(n24933), .op(n24649) );
  nor2_1 U24811 ( .ip1(n24648), .ip2(n24649), .op(n24907) );
  inv_1 U24812 ( .ip(n20743), .op(n20744) );
  nand2_1 U24813 ( .ip1(n20745), .ip2(n20744), .op(n20761) );
  inv_1 U24814 ( .ip(n20746), .op(n20748) );
  nor2_1 U24815 ( .ip1(n20748), .ip2(n20747), .op(n20753) );
  inv_1 U24816 ( .ip(n20749), .op(n20750) );
  nor2_1 U24817 ( .ip1(n20751), .ip2(n20750), .op(n20752) );
  not_ab_or_c_or_d U24818 ( .ip1(n20755), .ip2(n20754), .ip3(n20753), .ip4(
        n20752), .op(n20760) );
  nand3_1 U24819 ( .ip1(n20758), .ip2(n20757), .ip3(n20756), .op(n20759) );
  nand3_1 U24820 ( .ip1(n20761), .ip2(n20760), .ip3(n20759), .op(n24909) );
  nand2_1 U24821 ( .ip1(n24907), .ip2(n24909), .op(n24940) );
  nor2_1 U24822 ( .ip1(n24939), .ip2(n24940), .op(n24950) );
  nor2_1 U24823 ( .ip1(\x[73][14] ), .ip2(n23938), .op(n20762) );
  or2_1 U24824 ( .ip1(\x[73][15] ), .ip2(n20762), .op(n20764) );
  or2_1 U24825 ( .ip1(n23143), .ip2(n20762), .op(n20763) );
  nand2_1 U24826 ( .ip1(n20764), .ip2(n20763), .op(n20831) );
  nand2_1 U24827 ( .ip1(\x[73][14] ), .ip2(n24327), .op(n20825) );
  or2_1 U24828 ( .ip1(\x[73][13] ), .ip2(n24137), .op(n20767) );
  inv_1 U24829 ( .ip(\x[73][12] ), .op(n20765) );
  nand2_1 U24830 ( .ip1(n17845), .ip2(n20765), .op(n20766) );
  nand2_1 U24831 ( .ip1(n20767), .ip2(n20766), .op(n20827) );
  and2_1 U24832 ( .ip1(n24332), .ip2(\x[73][13] ), .op(n20805) );
  nand2_1 U24833 ( .ip1(\x[73][9] ), .ip2(n23981), .op(n20795) );
  nor2_1 U24834 ( .ip1(\x[73][9] ), .ip2(n24269), .op(n20790) );
  inv_1 U24835 ( .ip(\x[73][8] ), .op(n20768) );
  nor3_1 U24836 ( .ip1(sig_in[8]), .ip2(n20790), .ip3(n20768), .op(n20793) );
  and2_1 U24837 ( .ip1(n24461), .ip2(\x[73][7] ), .op(n20787) );
  inv_1 U24838 ( .ip(\x[73][5] ), .op(n20785) );
  nor2_1 U24839 ( .ip1(sig_in[5]), .ip2(n20785), .op(n20782) );
  inv_1 U24840 ( .ip(\x[73][3] ), .op(n20780) );
  and2_1 U24841 ( .ip1(n23659), .ip2(\x[73][2] ), .op(n20777) );
  inv_1 U24842 ( .ip(\x[73][1] ), .op(n20770) );
  inv_1 U24843 ( .ip(\x[73][0] ), .op(n20769) );
  not_ab_or_c_or_d U24844 ( .ip1(n24467), .ip2(n20770), .ip3(sig_in[0]), .ip4(
        n20769), .op(n20771) );
  or2_1 U24845 ( .ip1(\x[73][1] ), .ip2(n20771), .op(n20773) );
  or2_1 U24846 ( .ip1(n20652), .ip2(n20771), .op(n20772) );
  nand2_1 U24847 ( .ip1(n20773), .ip2(n20772), .op(n20775) );
  nor2_1 U24848 ( .ip1(\x[73][2] ), .ip2(n23717), .op(n20774) );
  nor2_1 U24849 ( .ip1(n20775), .ip2(n20774), .op(n20776) );
  not_ab_or_c_or_d U24850 ( .ip1(\x[73][3] ), .ip2(n22525), .ip3(n20777), 
        .ip4(n20776), .op(n20779) );
  nor2_1 U24851 ( .ip1(\x[73][4] ), .ip2(n24256), .op(n20778) );
  not_ab_or_c_or_d U24852 ( .ip1(n24251), .ip2(n20780), .ip3(n20779), .ip4(
        n20778), .op(n20781) );
  not_ab_or_c_or_d U24853 ( .ip1(\x[73][4] ), .ip2(n24347), .ip3(n20782), 
        .ip4(n20781), .op(n20784) );
  nor2_1 U24854 ( .ip1(\x[73][6] ), .ip2(n23509), .op(n20783) );
  not_ab_or_c_or_d U24855 ( .ip1(n22833), .ip2(n20785), .ip3(n20784), .ip4(
        n20783), .op(n20786) );
  not_ab_or_c_or_d U24856 ( .ip1(\x[73][6] ), .ip2(n24045), .ip3(n20787), 
        .ip4(n20786), .op(n20791) );
  nor2_1 U24857 ( .ip1(\x[73][8] ), .ip2(n24491), .op(n20789) );
  nor2_1 U24858 ( .ip1(\x[73][7] ), .ip2(n24492), .op(n20788) );
  nor4_1 U24859 ( .ip1(n20791), .ip2(n20790), .ip3(n20789), .ip4(n20788), .op(
        n20792) );
  not_ab_or_c_or_d U24860 ( .ip1(\x[73][10] ), .ip2(n20880), .ip3(n20793), 
        .ip4(n20792), .op(n20794) );
  nand2_1 U24861 ( .ip1(n20795), .ip2(n20794), .op(n20801) );
  nor2_1 U24862 ( .ip1(\x[73][10] ), .ip2(n24457), .op(n20796) );
  or2_1 U24863 ( .ip1(sig_in[11]), .ip2(n20796), .op(n20799) );
  inv_1 U24864 ( .ip(\x[73][11] ), .op(n20797) );
  or2_1 U24865 ( .ip1(n20797), .ip2(n20796), .op(n20798) );
  nand2_1 U24866 ( .ip1(n20799), .ip2(n20798), .op(n20800) );
  nand2_1 U24867 ( .ip1(n20801), .ip2(n20800), .op(n20803) );
  nand2_1 U24868 ( .ip1(\x[73][11] ), .ip2(n21793), .op(n20802) );
  nand2_1 U24869 ( .ip1(n20803), .ip2(n20802), .op(n20804) );
  not_ab_or_c_or_d U24870 ( .ip1(\x[73][12] ), .ip2(n24449), .ip3(n20805), 
        .ip4(n20804), .op(n20826) );
  or2_1 U24871 ( .ip1(n20827), .ip2(n20826), .op(n20806) );
  nand2_1 U24872 ( .ip1(n20825), .ip2(n20806), .op(n20811) );
  inv_1 U24873 ( .ip(n20807), .op(n20809) );
  nor2_1 U24874 ( .ip1(n20809), .ip2(n20808), .op(n20810) );
  nor2_1 U24875 ( .ip1(\x[73][15] ), .ip2(n24329), .op(n20830) );
  not_ab_or_c_or_d U24876 ( .ip1(n20831), .ip2(n20811), .ip3(n20810), .ip4(
        n20830), .op(n20819) );
  nand2_1 U24877 ( .ip1(n20813), .ip2(n20812), .op(n20815) );
  nand2_1 U24878 ( .ip1(n20815), .ip2(n20814), .op(n20817) );
  nand2_1 U24879 ( .ip1(n20817), .ip2(n20816), .op(n20818) );
  nand2_1 U24880 ( .ip1(n20819), .ip2(n20818), .op(n24952) );
  nand2_1 U24881 ( .ip1(n20821), .ip2(n20820), .op(n20823) );
  nand2_1 U24882 ( .ip1(n20823), .ip2(n20822), .op(n20840) );
  inv_1 U24883 ( .ip(n20830), .op(n20824) );
  nand2_1 U24884 ( .ip1(n20825), .ip2(n20824), .op(n20829) );
  nor2_1 U24885 ( .ip1(n20827), .ip2(n20826), .op(n20828) );
  nor2_1 U24886 ( .ip1(n20829), .ip2(n20828), .op(n20833) );
  nor2_1 U24887 ( .ip1(n20831), .ip2(n20830), .op(n20832) );
  nor2_1 U24888 ( .ip1(n20833), .ip2(n20832), .op(n20839) );
  inv_1 U24889 ( .ip(n20834), .op(n20835) );
  nand3_1 U24890 ( .ip1(n20837), .ip2(n20836), .ip3(n20835), .op(n20838) );
  nand3_1 U24891 ( .ip1(n20840), .ip2(n20839), .ip3(n20838), .op(n24951) );
  nand3_1 U24892 ( .ip1(n24950), .ip2(n24952), .ip3(n24951), .op(n24949) );
  nor2_1 U24893 ( .ip1(n24947), .ip2(n24949), .op(n27567) );
  inv_1 U24894 ( .ip(n20841), .op(n20900) );
  inv_1 U24895 ( .ip(n20842), .op(n20899) );
  and3_1 U24896 ( .ip1(n20845), .ip2(n20844), .ip3(n20843), .op(n20898) );
  nand2_1 U24897 ( .ip1(n24332), .ip2(\x[86][13] ), .op(n20847) );
  nand2_1 U24898 ( .ip1(\x[86][12] ), .ip2(n24233), .op(n20846) );
  nand2_1 U24899 ( .ip1(n20847), .ip2(n20846), .op(n21615) );
  nand2_1 U24900 ( .ip1(\x[86][11] ), .ip2(n21793), .op(n20849) );
  nand2_1 U24901 ( .ip1(\x[86][10] ), .ip2(n23146), .op(n20848) );
  nand2_1 U24902 ( .ip1(n20849), .ip2(n20848), .op(n20879) );
  and2_1 U24903 ( .ip1(n24335), .ip2(\x[86][2] ), .op(n20858) );
  inv_1 U24904 ( .ip(\x[86][1] ), .op(n20851) );
  inv_1 U24905 ( .ip(\x[86][0] ), .op(n20850) );
  not_ab_or_c_or_d U24906 ( .ip1(n24467), .ip2(n20851), .ip3(n23195), .ip4(
        n20850), .op(n20852) );
  or2_1 U24907 ( .ip1(\x[86][1] ), .ip2(n20852), .op(n20854) );
  or2_1 U24908 ( .ip1(n20652), .ip2(n20852), .op(n20853) );
  nand2_1 U24909 ( .ip1(n20854), .ip2(n20853), .op(n20856) );
  nor2_1 U24910 ( .ip1(\x[86][2] ), .ip2(n23717), .op(n20855) );
  nor2_1 U24911 ( .ip1(n20856), .ip2(n20855), .op(n20857) );
  not_ab_or_c_or_d U24912 ( .ip1(\x[86][3] ), .ip2(n24476), .ip3(n20858), 
        .ip4(n20857), .op(n20861) );
  nor2_1 U24913 ( .ip1(\x[86][5] ), .ip2(n24119), .op(n20862) );
  nor2_1 U24914 ( .ip1(\x[86][3] ), .ip2(n24342), .op(n20860) );
  nor2_1 U24915 ( .ip1(\x[86][4] ), .ip2(n23860), .op(n20859) );
  nor4_1 U24916 ( .ip1(n20861), .ip2(n20862), .ip3(n20860), .ip4(n20859), .op(
        n20868) );
  nand2_1 U24917 ( .ip1(n23600), .ip2(\x[86][5] ), .op(n20866) );
  inv_1 U24918 ( .ip(n20862), .op(n20863) );
  nand3_1 U24919 ( .ip1(\x[86][4] ), .ip2(n23721), .ip3(n20863), .op(n20865)
         );
  nand2_1 U24920 ( .ip1(\x[86][7] ), .ip2(n24044), .op(n20864) );
  nand3_1 U24921 ( .ip1(n20866), .ip2(n20865), .ip3(n20864), .op(n20867) );
  not_ab_or_c_or_d U24922 ( .ip1(\x[86][6] ), .ip2(n24045), .ip3(n20868), 
        .ip4(n20867), .op(n20872) );
  not_ab_or_c_or_d U24923 ( .ip1(\x[86][7] ), .ip2(n24044), .ip3(\x[86][6] ), 
        .ip4(n23509), .op(n20871) );
  nor2_1 U24924 ( .ip1(\x[86][7] ), .ip2(n24492), .op(n20870) );
  nor2_1 U24925 ( .ip1(\x[86][8] ), .ip2(n24491), .op(n20869) );
  or4_1 U24926 ( .ip1(n20872), .ip2(n20871), .ip3(n20870), .ip4(n20869), .op(
        n20873) );
  nor2_1 U24927 ( .ip1(\x[86][9] ), .ip2(n24164), .op(n20874) );
  or2_1 U24928 ( .ip1(n20873), .ip2(n20874), .op(n20877) );
  nand2_1 U24929 ( .ip1(\x[86][8] ), .ip2(n24491), .op(n20875) );
  or2_1 U24930 ( .ip1(n20875), .ip2(n20874), .op(n20876) );
  nand2_1 U24931 ( .ip1(n20877), .ip2(n20876), .op(n20878) );
  not_ab_or_c_or_d U24932 ( .ip1(\x[86][9] ), .ip2(n24043), .ip3(n20879), 
        .ip4(n20878), .op(n20884) );
  nor2_1 U24933 ( .ip1(n24456), .ip2(\x[86][11] ), .op(n20882) );
  not_ab_or_c_or_d U24934 ( .ip1(\x[86][11] ), .ip2(n24136), .ip3(\x[86][10] ), 
        .ip4(n20880), .op(n20881) );
  or2_1 U24935 ( .ip1(n20882), .ip2(n20881), .op(n20883) );
  nor2_1 U24936 ( .ip1(n20884), .ip2(n20883), .op(n21618) );
  or2_1 U24937 ( .ip1(n21615), .ip2(n21618), .op(n20889) );
  nor2_1 U24938 ( .ip1(\x[86][13] ), .ip2(n24376), .op(n20885) );
  or2_1 U24939 ( .ip1(n17845), .ip2(n20885), .op(n20888) );
  inv_1 U24940 ( .ip(\x[86][12] ), .op(n20886) );
  or2_1 U24941 ( .ip1(n20886), .ip2(n20885), .op(n20887) );
  nand2_1 U24942 ( .ip1(n20888), .ip2(n20887), .op(n21617) );
  nand2_1 U24943 ( .ip1(n20889), .ip2(n21617), .op(n20892) );
  nor2_1 U24944 ( .ip1(\x[86][15] ), .ip2(n24180), .op(n20894) );
  or2_1 U24945 ( .ip1(\x[86][14] ), .ip2(n20894), .op(n20891) );
  or2_1 U24946 ( .ip1(n24185), .ip2(n20894), .op(n20890) );
  nand2_1 U24947 ( .ip1(n20891), .ip2(n20890), .op(n21621) );
  nand2_1 U24948 ( .ip1(n20892), .ip2(n21621), .op(n20896) );
  nand2_1 U24949 ( .ip1(\x[86][15] ), .ip2(n24186), .op(n21623) );
  or2_1 U24950 ( .ip1(n24185), .ip2(\x[86][14] ), .op(n20893) );
  and2_1 U24951 ( .ip1(n21623), .ip2(n20893), .op(n21616) );
  or2_1 U24952 ( .ip1(n21616), .ip2(n20894), .op(n20895) );
  nand2_1 U24953 ( .ip1(n20896), .ip2(n20895), .op(n20897) );
  not_ab_or_c_or_d U24954 ( .ip1(n20900), .ip2(n20899), .ip3(n20898), .ip4(
        n20897), .op(n24569) );
  nor2_1 U24955 ( .ip1(\x[88][13] ), .ip2(n24137), .op(n20901) );
  or2_1 U24956 ( .ip1(n17845), .ip2(n20901), .op(n20904) );
  inv_1 U24957 ( .ip(\x[88][12] ), .op(n20902) );
  or2_1 U24958 ( .ip1(n20902), .ip2(n20901), .op(n20903) );
  nand2_1 U24959 ( .ip1(n20904), .ip2(n20903), .op(n21596) );
  inv_1 U24960 ( .ip(\x[88][11] ), .op(n20931) );
  and2_1 U24961 ( .ip1(n24451), .ip2(\x[88][10] ), .op(n20928) );
  inv_1 U24962 ( .ip(\x[88][9] ), .op(n20926) );
  and2_1 U24963 ( .ip1(n23804), .ip2(\x[88][8] ), .op(n20923) );
  nor2_1 U24964 ( .ip1(\x[88][5] ), .ip2(n23283), .op(n20914) );
  inv_1 U24965 ( .ip(\x[88][4] ), .op(n20905) );
  nor3_1 U24966 ( .ip1(n24462), .ip2(n20914), .ip3(n20905), .op(n20917) );
  and2_1 U24967 ( .ip1(n23659), .ip2(\x[88][2] ), .op(n20911) );
  nand2_1 U24968 ( .ip1(\x[88][1] ), .ip2(n20652), .op(n20909) );
  nand2_1 U24969 ( .ip1(\x[88][0] ), .ip2(n24143), .op(n20908) );
  nor2_1 U24970 ( .ip1(\x[88][2] ), .ip2(n23717), .op(n20907) );
  nor2_1 U24971 ( .ip1(\x[88][1] ), .ip2(n20652), .op(n20906) );
  not_ab_or_c_or_d U24972 ( .ip1(n20909), .ip2(n20908), .ip3(n20907), .ip4(
        n20906), .op(n20910) );
  not_ab_or_c_or_d U24973 ( .ip1(\x[88][3] ), .ip2(n22525), .ip3(n20911), 
        .ip4(n20910), .op(n20915) );
  nor2_1 U24974 ( .ip1(\x[88][3] ), .ip2(n24342), .op(n20913) );
  nor2_1 U24975 ( .ip1(\x[88][4] ), .ip2(n24347), .op(n20912) );
  nor4_1 U24976 ( .ip1(n20915), .ip2(n20914), .ip3(n20913), .ip4(n20912), .op(
        n20916) );
  not_ab_or_c_or_d U24977 ( .ip1(\x[88][6] ), .ip2(n24045), .ip3(n20917), 
        .ip4(n20916), .op(n20921) );
  nand2_1 U24978 ( .ip1(\x[88][5] ), .ip2(n24119), .op(n20920) );
  nor2_1 U24979 ( .ip1(\x[88][7] ), .ip2(n24044), .op(n20919) );
  nor2_1 U24980 ( .ip1(\x[88][6] ), .ip2(n23509), .op(n20918) );
  not_ab_or_c_or_d U24981 ( .ip1(n20921), .ip2(n20920), .ip3(n20919), .ip4(
        n20918), .op(n20922) );
  not_ab_or_c_or_d U24982 ( .ip1(\x[88][7] ), .ip2(n24142), .ip3(n20923), 
        .ip4(n20922), .op(n20925) );
  nor2_1 U24983 ( .ip1(\x[88][8] ), .ip2(n24491), .op(n20924) );
  not_ab_or_c_or_d U24984 ( .ip1(sig_in[9]), .ip2(n20926), .ip3(n20925), .ip4(
        n20924), .op(n20927) );
  not_ab_or_c_or_d U24985 ( .ip1(\x[88][9] ), .ip2(n24269), .ip3(n20928), 
        .ip4(n20927), .op(n20930) );
  nor2_1 U24986 ( .ip1(\x[88][10] ), .ip2(n24457), .op(n20929) );
  not_ab_or_c_or_d U24987 ( .ip1(sig_in[11]), .ip2(n20931), .ip3(n20930), 
        .ip4(n20929), .op(n20932) );
  or2_1 U24988 ( .ip1(\x[88][11] ), .ip2(n20932), .op(n20934) );
  or2_1 U24989 ( .ip1(n24136), .ip2(n20932), .op(n20933) );
  nand2_1 U24990 ( .ip1(n20934), .ip2(n20933), .op(n21594) );
  nand2_1 U24991 ( .ip1(\x[88][12] ), .ip2(n24450), .op(n21602) );
  nand2_1 U24992 ( .ip1(n21594), .ip2(n21602), .op(n20937) );
  nor2_1 U24993 ( .ip1(\x[88][15] ), .ip2(n24180), .op(n21590) );
  nand2_1 U24994 ( .ip1(\x[88][14] ), .ip2(n24230), .op(n20936) );
  nand2_1 U24995 ( .ip1(\x[88][13] ), .ip2(n24235), .op(n20935) );
  nand2_1 U24996 ( .ip1(n20936), .ip2(n20935), .op(n21601) );
  not_ab_or_c_or_d U24997 ( .ip1(n21596), .ip2(n20937), .ip3(n21590), .ip4(
        n21601), .op(n20994) );
  nand2_1 U24998 ( .ip1(n23143), .ip2(\x[88][15] ), .op(n21605) );
  inv_1 U24999 ( .ip(n21605), .op(n20938) );
  or2_1 U25000 ( .ip1(sig_in[14]), .ip2(n20938), .op(n20941) );
  inv_1 U25001 ( .ip(\x[88][14] ), .op(n20939) );
  or2_1 U25002 ( .ip1(n20939), .ip2(n20938), .op(n20940) );
  nand2_1 U25003 ( .ip1(n20941), .ip2(n20940), .op(n21597) );
  nor2_1 U25004 ( .ip1(n21597), .ip2(n21590), .op(n20993) );
  nand2_1 U25005 ( .ip1(n24327), .ip2(\x[87][14] ), .op(n20944) );
  nor2_1 U25006 ( .ip1(n24384), .ip2(\x[87][15] ), .op(n20950) );
  inv_1 U25007 ( .ip(n20950), .op(n20943) );
  nand2_1 U25008 ( .ip1(\x[87][13] ), .ip2(n24081), .op(n20942) );
  nand3_1 U25009 ( .ip1(n20944), .ip2(n20943), .ip3(n20942), .op(n21620) );
  or2_1 U25010 ( .ip1(\x[87][12] ), .ip2(n21620), .op(n20946) );
  or2_1 U25011 ( .ip1(n24449), .ip2(n21620), .op(n20945) );
  nand2_1 U25012 ( .ip1(n20946), .ip2(n20945), .op(n21610) );
  nor2_1 U25013 ( .ip1(\x[87][14] ), .ip2(n23938), .op(n20947) );
  or2_1 U25014 ( .ip1(\x[87][15] ), .ip2(n20947), .op(n20949) );
  or2_1 U25015 ( .ip1(n24329), .ip2(n20947), .op(n20948) );
  nand2_1 U25016 ( .ip1(n20949), .ip2(n20948), .op(n20990) );
  nor2_1 U25017 ( .ip1(n20950), .ip2(n20990), .op(n21614) );
  nor2_1 U25018 ( .ip1(n21610), .ip2(n21614), .op(n20992) );
  nand2_1 U25019 ( .ip1(\x[87][10] ), .ip2(n23146), .op(n20952) );
  nand2_1 U25020 ( .ip1(\x[87][11] ), .ip2(n21793), .op(n20951) );
  nand2_1 U25021 ( .ip1(n20952), .ip2(n20951), .op(n20977) );
  nor3_1 U25022 ( .ip1(\x[87][9] ), .ip2(n24455), .ip3(n20977), .op(n20985) );
  not_ab_or_c_or_d U25023 ( .ip1(\x[87][11] ), .ip2(n24136), .ip3(\x[87][10] ), 
        .ip4(n24370), .op(n20984) );
  nor2_1 U25024 ( .ip1(\x[87][11] ), .ip2(n24239), .op(n20983) );
  inv_1 U25025 ( .ip(\x[87][5] ), .op(n20967) );
  nor2_1 U25026 ( .ip1(sig_in[5]), .ip2(n20967), .op(n20964) );
  nor2_1 U25027 ( .ip1(\x[87][4] ), .ip2(n23721), .op(n20962) );
  not_ab_or_c_or_d U25028 ( .ip1(\x[87][3] ), .ip2(n24476), .ip3(\x[87][2] ), 
        .ip4(n24470), .op(n20961) );
  nor2_1 U25029 ( .ip1(\x[87][3] ), .ip2(n24342), .op(n20960) );
  inv_1 U25030 ( .ip(\x[87][1] ), .op(n20954) );
  inv_1 U25031 ( .ip(\x[87][0] ), .op(n20953) );
  not_ab_or_c_or_d U25032 ( .ip1(n24467), .ip2(n20954), .ip3(n23195), .ip4(
        n20953), .op(n20958) );
  nand2_1 U25033 ( .ip1(\x[87][3] ), .ip2(n22795), .op(n20956) );
  nand2_1 U25034 ( .ip1(\x[87][1] ), .ip2(n21685), .op(n20955) );
  nand2_1 U25035 ( .ip1(n20956), .ip2(n20955), .op(n20957) );
  not_ab_or_c_or_d U25036 ( .ip1(\x[87][2] ), .ip2(n24107), .ip3(n20958), 
        .ip4(n20957), .op(n20959) );
  nor4_1 U25037 ( .ip1(n20962), .ip2(n20961), .ip3(n20960), .ip4(n20959), .op(
        n20963) );
  not_ab_or_c_or_d U25038 ( .ip1(\x[87][4] ), .ip2(n23860), .ip3(n20964), 
        .ip4(n20963), .op(n20966) );
  nor2_1 U25039 ( .ip1(\x[87][6] ), .ip2(n23509), .op(n20965) );
  not_ab_or_c_or_d U25040 ( .ip1(sig_in[5]), .ip2(n20967), .ip3(n20966), .ip4(
        n20965), .op(n20968) );
  or2_1 U25041 ( .ip1(\x[87][6] ), .ip2(n20968), .op(n20970) );
  or2_1 U25042 ( .ip1(n24045), .ip2(n20968), .op(n20969) );
  nand2_1 U25043 ( .ip1(n20970), .ip2(n20969), .op(n20972) );
  nor2_1 U25044 ( .ip1(\x[87][7] ), .ip2(n24492), .op(n20971) );
  nor2_1 U25045 ( .ip1(n20972), .ip2(n20971), .op(n20974) );
  and2_1 U25046 ( .ip1(n23804), .ip2(\x[87][8] ), .op(n20973) );
  not_ab_or_c_or_d U25047 ( .ip1(\x[87][7] ), .ip2(n24142), .ip3(n20974), 
        .ip4(n20973), .op(n20976) );
  nor2_1 U25048 ( .ip1(n24358), .ip2(\x[87][8] ), .op(n20975) );
  nor2_1 U25049 ( .ip1(n20976), .ip2(n20975), .op(n20981) );
  inv_1 U25050 ( .ip(n20977), .op(n20979) );
  nand2_1 U25051 ( .ip1(\x[87][9] ), .ip2(n24164), .op(n20978) );
  nand2_1 U25052 ( .ip1(n20979), .ip2(n20978), .op(n20980) );
  nor2_1 U25053 ( .ip1(n20981), .ip2(n20980), .op(n20982) );
  nor4_1 U25054 ( .ip1(n20985), .ip2(n20984), .ip3(n20983), .ip4(n20982), .op(
        n21612) );
  nor2_1 U25055 ( .ip1(\x[87][13] ), .ip2(n24137), .op(n20986) );
  or2_1 U25056 ( .ip1(n17845), .ip2(n20986), .op(n20989) );
  inv_1 U25057 ( .ip(\x[87][12] ), .op(n20987) );
  or2_1 U25058 ( .ip1(n20987), .ip2(n20986), .op(n20988) );
  nand2_1 U25059 ( .ip1(n20989), .ip2(n20988), .op(n21619) );
  and3_1 U25060 ( .ip1(n20990), .ip2(n21612), .ip3(n21619), .op(n20991) );
  nor4_1 U25061 ( .ip1(n20994), .ip2(n20993), .ip3(n20992), .ip4(n20991), .op(
        n24526) );
  and2_1 U25062 ( .ip1(n24332), .ip2(\x[90][13] ), .op(n20995) );
  nor2_1 U25063 ( .ip1(\x[90][15] ), .ip2(n24180), .op(n21001) );
  not_ab_or_c_or_d U25064 ( .ip1(\x[90][14] ), .ip2(n24382), .ip3(n20995), 
        .ip4(n21001), .op(n21092) );
  nor2_1 U25065 ( .ip1(\x[90][13] ), .ip2(n24376), .op(n20997) );
  nor2_1 U25066 ( .ip1(\x[90][12] ), .ip2(n24079), .op(n20996) );
  nor2_1 U25067 ( .ip1(n20997), .ip2(n20996), .op(n21585) );
  inv_1 U25068 ( .ip(n21585), .op(n21091) );
  and2_1 U25069 ( .ip1(n24186), .ip2(\x[90][15] ), .op(n21568) );
  or2_1 U25070 ( .ip1(sig_in[14]), .ip2(n21568), .op(n21000) );
  inv_1 U25071 ( .ip(\x[90][14] ), .op(n20998) );
  or2_1 U25072 ( .ip1(n20998), .ip2(n21568), .op(n20999) );
  nand2_1 U25073 ( .ip1(n21000), .ip2(n20999), .op(n21584) );
  nor2_1 U25074 ( .ip1(n21001), .ip2(n21584), .op(n21090) );
  inv_1 U25075 ( .ip(n21092), .op(n21002) );
  or2_1 U25076 ( .ip1(\x[90][12] ), .ip2(n21002), .op(n21004) );
  or2_1 U25077 ( .ip1(n24449), .ip2(n21002), .op(n21003) );
  nand2_1 U25078 ( .ip1(n21004), .ip2(n21003), .op(n21567) );
  inv_1 U25079 ( .ip(\x[90][11] ), .op(n21038) );
  and2_1 U25080 ( .ip1(n24451), .ip2(\x[90][10] ), .op(n21035) );
  inv_1 U25081 ( .ip(\x[90][9] ), .op(n21033) );
  inv_1 U25082 ( .ip(\x[90][7] ), .op(n21025) );
  nor2_1 U25083 ( .ip1(n17732), .ip2(n21025), .op(n21023) );
  inv_1 U25084 ( .ip(\x[90][5] ), .op(n21021) );
  nor2_1 U25085 ( .ip1(sig_in[5]), .ip2(n21021), .op(n21018) );
  inv_1 U25086 ( .ip(\x[90][3] ), .op(n21016) );
  inv_1 U25087 ( .ip(\x[90][1] ), .op(n21006) );
  nor2_1 U25088 ( .ip1(n24464), .ip2(n21006), .op(n21008) );
  inv_1 U25089 ( .ip(\x[90][0] ), .op(n21005) );
  not_ab_or_c_or_d U25090 ( .ip1(n24467), .ip2(n21006), .ip3(sig_in[0]), .ip4(
        n21005), .op(n21007) );
  not_ab_or_c_or_d U25091 ( .ip1(\x[90][2] ), .ip2(n24107), .ip3(n21008), 
        .ip4(n21007), .op(n21010) );
  nor2_1 U25092 ( .ip1(\x[90][2] ), .ip2(n23717), .op(n21009) );
  nor2_1 U25093 ( .ip1(n21010), .ip2(n21009), .op(n21011) );
  or2_1 U25094 ( .ip1(\x[90][3] ), .ip2(n21011), .op(n21013) );
  or2_1 U25095 ( .ip1(n24476), .ip2(n21011), .op(n21012) );
  nand2_1 U25096 ( .ip1(n21013), .ip2(n21012), .op(n21015) );
  nor2_1 U25097 ( .ip1(\x[90][4] ), .ip2(n24256), .op(n21014) );
  not_ab_or_c_or_d U25098 ( .ip1(n23251), .ip2(n21016), .ip3(n21015), .ip4(
        n21014), .op(n21017) );
  not_ab_or_c_or_d U25099 ( .ip1(\x[90][4] ), .ip2(n24347), .ip3(n21018), 
        .ip4(n21017), .op(n21020) );
  nor2_1 U25100 ( .ip1(\x[90][6] ), .ip2(n23509), .op(n21019) );
  not_ab_or_c_or_d U25101 ( .ip1(n22833), .ip2(n21021), .ip3(n21020), .ip4(
        n21019), .op(n21022) );
  not_ab_or_c_or_d U25102 ( .ip1(\x[90][6] ), .ip2(n24045), .ip3(n21023), 
        .ip4(n21022), .op(n21024) );
  or2_1 U25103 ( .ip1(n17732), .ip2(n21024), .op(n21027) );
  or2_1 U25104 ( .ip1(n21025), .ip2(n21024), .op(n21026) );
  nand2_1 U25105 ( .ip1(n21027), .ip2(n21026), .op(n21028) );
  or2_1 U25106 ( .ip1(\x[90][8] ), .ip2(n21028), .op(n21030) );
  or2_1 U25107 ( .ip1(n24100), .ip2(n21028), .op(n21029) );
  nand2_1 U25108 ( .ip1(n21030), .ip2(n21029), .op(n21032) );
  nor2_1 U25109 ( .ip1(\x[90][8] ), .ip2(n24491), .op(n21031) );
  not_ab_or_c_or_d U25110 ( .ip1(sig_in[9]), .ip2(n21033), .ip3(n21032), .ip4(
        n21031), .op(n21034) );
  not_ab_or_c_or_d U25111 ( .ip1(\x[90][9] ), .ip2(n24269), .ip3(n21035), 
        .ip4(n21034), .op(n21037) );
  nor2_1 U25112 ( .ip1(\x[90][10] ), .ip2(n24457), .op(n21036) );
  not_ab_or_c_or_d U25113 ( .ip1(sig_in[11]), .ip2(n21038), .ip3(n21037), 
        .ip4(n21036), .op(n21039) );
  or2_1 U25114 ( .ip1(\x[90][11] ), .ip2(n21039), .op(n21041) );
  or2_1 U25115 ( .ip1(n24136), .ip2(n21039), .op(n21040) );
  nand2_1 U25116 ( .ip1(n21041), .ip2(n21040), .op(n21582) );
  nand2_1 U25117 ( .ip1(n21567), .ip2(n21582), .op(n21088) );
  nor2_1 U25118 ( .ip1(\x[89][13] ), .ip2(n24376), .op(n21042) );
  or2_1 U25119 ( .ip1(sig_in[12]), .ip2(n21042), .op(n21045) );
  inv_1 U25120 ( .ip(\x[89][12] ), .op(n21043) );
  or2_1 U25121 ( .ip1(n21043), .ip2(n21042), .op(n21044) );
  nand2_1 U25122 ( .ip1(n21045), .ip2(n21044), .op(n21598) );
  nor2_1 U25123 ( .ip1(\x[89][14] ), .ip2(n23938), .op(n21046) );
  or2_1 U25124 ( .ip1(\x[89][15] ), .ip2(n21046), .op(n21048) );
  or2_1 U25125 ( .ip1(n24180), .ip2(n21046), .op(n21047) );
  nand2_1 U25126 ( .ip1(n21048), .ip2(n21047), .op(n21085) );
  nand2_1 U25127 ( .ip1(\x[89][10] ), .ip2(n23146), .op(n21077) );
  nand2_1 U25128 ( .ip1(n21077), .ip2(n17981), .op(n21080) );
  and2_1 U25129 ( .ip1(n23804), .ip2(\x[89][8] ), .op(n21071) );
  inv_1 U25130 ( .ip(\x[89][7] ), .op(n21068) );
  nor2_1 U25131 ( .ip1(n17732), .ip2(n21068), .op(n21065) );
  inv_1 U25132 ( .ip(\x[89][3] ), .op(n21055) );
  nor2_1 U25133 ( .ip1(\x[89][2] ), .ip2(n23717), .op(n21054) );
  inv_1 U25134 ( .ip(\x[89][1] ), .op(n21050) );
  nor2_1 U25135 ( .ip1(n24464), .ip2(n21050), .op(n21052) );
  inv_1 U25136 ( .ip(\x[89][0] ), .op(n21049) );
  not_ab_or_c_or_d U25137 ( .ip1(n24467), .ip2(n21050), .ip3(n23195), .ip4(
        n21049), .op(n21051) );
  not_ab_or_c_or_d U25138 ( .ip1(\x[89][2] ), .ip2(n24470), .ip3(n21052), 
        .ip4(n21051), .op(n21053) );
  not_ab_or_c_or_d U25139 ( .ip1(sig_in[3]), .ip2(n21055), .ip3(n21054), .ip4(
        n21053), .op(n21059) );
  nand2_1 U25140 ( .ip1(\x[89][5] ), .ip2(n24119), .op(n21057) );
  nand2_1 U25141 ( .ip1(\x[89][4] ), .ip2(n24256), .op(n21056) );
  nand2_1 U25142 ( .ip1(n21057), .ip2(n21056), .op(n21058) );
  not_ab_or_c_or_d U25143 ( .ip1(\x[89][3] ), .ip2(n22525), .ip3(n21059), 
        .ip4(n21058), .op(n21063) );
  nor2_1 U25144 ( .ip1(\x[89][5] ), .ip2(n23283), .op(n21062) );
  nor2_1 U25145 ( .ip1(\x[89][6] ), .ip2(n23770), .op(n21061) );
  not_ab_or_c_or_d U25146 ( .ip1(\x[89][5] ), .ip2(n24482), .ip3(\x[89][4] ), 
        .ip4(n24256), .op(n21060) );
  nor4_1 U25147 ( .ip1(n21063), .ip2(n21062), .ip3(n21061), .ip4(n21060), .op(
        n21064) );
  not_ab_or_c_or_d U25148 ( .ip1(\x[89][6] ), .ip2(n24045), .ip3(n21065), 
        .ip4(n21064), .op(n21067) );
  nor2_1 U25149 ( .ip1(\x[89][8] ), .ip2(n24491), .op(n21066) );
  not_ab_or_c_or_d U25150 ( .ip1(n17732), .ip2(n21068), .ip3(n21067), .ip4(
        n21066), .op(n21070) );
  inv_1 U25151 ( .ip(\x[89][9] ), .op(n21074) );
  nor2_1 U25152 ( .ip1(n21171), .ip2(n21074), .op(n21069) );
  nor3_1 U25153 ( .ip1(n21071), .ip2(n21070), .ip3(n21069), .op(n21076) );
  nor2_1 U25154 ( .ip1(\x[89][11] ), .ip2(n24371), .op(n21073) );
  nor2_1 U25155 ( .ip1(\x[89][10] ), .ip2(n24457), .op(n21072) );
  ab_or_c_or_d U25156 ( .ip1(n21171), .ip2(n21074), .ip3(n21073), .ip4(n21072), 
        .op(n21075) );
  nor2_1 U25157 ( .ip1(n21076), .ip2(n21075), .op(n21079) );
  nor2_1 U25158 ( .ip1(n21077), .ip2(n17981), .op(n21078) );
  not_ab_or_c_or_d U25159 ( .ip1(\x[89][11] ), .ip2(n21080), .ip3(n21079), 
        .ip4(n21078), .op(n21592) );
  inv_1 U25160 ( .ip(n21592), .op(n21081) );
  nand3_1 U25161 ( .ip1(n21598), .ip2(n21085), .ip3(n21081), .op(n21087) );
  and2_1 U25162 ( .ip1(n23895), .ip2(\x[89][13] ), .op(n21082) );
  nor2_1 U25163 ( .ip1(\x[89][15] ), .ip2(n24329), .op(n21084) );
  not_ab_or_c_or_d U25164 ( .ip1(\x[89][14] ), .ip2(n24382), .ip3(n21082), 
        .ip4(n21084), .op(n21600) );
  nand2_1 U25165 ( .ip1(\x[89][12] ), .ip2(n24450), .op(n21083) );
  and2_1 U25166 ( .ip1(n21600), .ip2(n21083), .op(n21593) );
  nor2_1 U25167 ( .ip1(n21085), .ip2(n21084), .op(n21591) );
  or2_1 U25168 ( .ip1(n21593), .ip2(n21591), .op(n21086) );
  nand3_1 U25169 ( .ip1(n21088), .ip2(n21087), .ip3(n21086), .op(n21089) );
  not_ab_or_c_or_d U25170 ( .ip1(n21092), .ip2(n21091), .ip3(n21090), .ip4(
        n21089), .op(n24556) );
  nand2_1 U25171 ( .ip1(\x[91][15] ), .ip2(n24186), .op(n21186) );
  and2_1 U25172 ( .ip1(n24332), .ip2(\x[91][13] ), .op(n21093) );
  nor2_1 U25173 ( .ip1(\x[91][15] ), .ip2(n24180), .op(n21564) );
  not_ab_or_c_or_d U25174 ( .ip1(\x[91][14] ), .ip2(n24382), .ip3(n21093), 
        .ip4(n21564), .op(n21579) );
  nand2_1 U25175 ( .ip1(\x[91][12] ), .ip2(n24079), .op(n21578) );
  nand2_1 U25176 ( .ip1(n21579), .ip2(n21578), .op(n21185) );
  inv_1 U25177 ( .ip(\x[91][11] ), .op(n21097) );
  nor2_1 U25178 ( .ip1(n17981), .ip2(n21097), .op(n21100) );
  or2_1 U25179 ( .ip1(\x[91][10] ), .ip2(n21100), .op(n21095) );
  or2_1 U25180 ( .ip1(n23980), .ip2(n21100), .op(n21094) );
  nand2_1 U25181 ( .ip1(n21095), .ip2(n21094), .op(n21104) );
  nor2_1 U25182 ( .ip1(\x[91][9] ), .ip2(n24269), .op(n21129) );
  nor2_1 U25183 ( .ip1(\x[91][10] ), .ip2(n24457), .op(n21096) );
  or2_1 U25184 ( .ip1(sig_in[11]), .ip2(n21096), .op(n21099) );
  or2_1 U25185 ( .ip1(n21097), .ip2(n21096), .op(n21098) );
  nand2_1 U25186 ( .ip1(n21099), .ip2(n21098), .op(n21130) );
  nor2_1 U25187 ( .ip1(n21100), .ip2(n21130), .op(n21572) );
  nand2_1 U25188 ( .ip1(\x[91][9] ), .ip2(n24043), .op(n21101) );
  nand2_1 U25189 ( .ip1(n21104), .ip2(n21101), .op(n21569) );
  or2_1 U25190 ( .ip1(\x[91][8] ), .ip2(n21569), .op(n21103) );
  or2_1 U25191 ( .ip1(n24100), .ip2(n21569), .op(n21102) );
  nand2_1 U25192 ( .ip1(n21103), .ip2(n21102), .op(n21574) );
  not_ab_or_c_or_d U25193 ( .ip1(n21104), .ip2(n21129), .ip3(n21572), .ip4(
        n21574), .op(n21133) );
  nor2_1 U25194 ( .ip1(\x[91][5] ), .ip2(n23283), .op(n21116) );
  inv_1 U25195 ( .ip(\x[91][4] ), .op(n21105) );
  nor3_1 U25196 ( .ip1(n24462), .ip2(n21116), .ip3(n21105), .op(n21120) );
  nor2_1 U25197 ( .ip1(\x[91][4] ), .ip2(n23860), .op(n21118) );
  nor2_1 U25198 ( .ip1(\x[91][3] ), .ip2(n24342), .op(n21117) );
  inv_1 U25199 ( .ip(\x[91][1] ), .op(n21107) );
  nor2_1 U25200 ( .ip1(n24464), .ip2(n21107), .op(n21109) );
  inv_1 U25201 ( .ip(\x[91][0] ), .op(n21106) );
  not_ab_or_c_or_d U25202 ( .ip1(n24467), .ip2(n21107), .ip3(n23195), .ip4(
        n21106), .op(n21108) );
  not_ab_or_c_or_d U25203 ( .ip1(\x[91][2] ), .ip2(n24470), .ip3(n21109), 
        .ip4(n21108), .op(n21111) );
  nor2_1 U25204 ( .ip1(\x[91][2] ), .ip2(n23717), .op(n21110) );
  nor2_1 U25205 ( .ip1(n21111), .ip2(n21110), .op(n21112) );
  or2_1 U25206 ( .ip1(\x[91][3] ), .ip2(n21112), .op(n21114) );
  or2_1 U25207 ( .ip1(n24476), .ip2(n21112), .op(n21113) );
  nand2_1 U25208 ( .ip1(n21114), .ip2(n21113), .op(n21115) );
  nor4_1 U25209 ( .ip1(n21118), .ip2(n21117), .ip3(n21116), .ip4(n21115), .op(
        n21119) );
  not_ab_or_c_or_d U25210 ( .ip1(\x[91][5] ), .ip2(n24482), .ip3(n21120), 
        .ip4(n21119), .op(n21124) );
  nand2_1 U25211 ( .ip1(\x[91][6] ), .ip2(n24485), .op(n21123) );
  nor2_1 U25212 ( .ip1(\x[91][6] ), .ip2(n23770), .op(n21122) );
  nor2_1 U25213 ( .ip1(\x[91][7] ), .ip2(n24492), .op(n21121) );
  not_ab_or_c_or_d U25214 ( .ip1(n21124), .ip2(n21123), .ip3(n21122), .ip4(
        n21121), .op(n21125) );
  or2_1 U25215 ( .ip1(\x[91][7] ), .ip2(n21125), .op(n21127) );
  or2_1 U25216 ( .ip1(n24142), .ip2(n21125), .op(n21126) );
  nand2_1 U25217 ( .ip1(n21127), .ip2(n21126), .op(n21573) );
  inv_1 U25218 ( .ip(n21573), .op(n21131) );
  nor2_1 U25219 ( .ip1(\x[91][8] ), .ip2(n24491), .op(n21128) );
  nor2_1 U25220 ( .ip1(n21129), .ip2(n21128), .op(n21570) );
  and3_1 U25221 ( .ip1(n21131), .ip2(n21130), .ip3(n21570), .op(n21132) );
  nor2_1 U25222 ( .ip1(n21133), .ip2(n21132), .op(n21137) );
  nor2_1 U25223 ( .ip1(\x[91][13] ), .ip2(n24137), .op(n21135) );
  nor2_1 U25224 ( .ip1(\x[91][12] ), .ip2(n24449), .op(n21134) );
  nor2_1 U25225 ( .ip1(n21135), .ip2(n21134), .op(n21575) );
  inv_1 U25226 ( .ip(n21575), .op(n21577) );
  or2_1 U25227 ( .ip1(n24382), .ip2(\x[91][14] ), .op(n21136) );
  nand2_1 U25228 ( .ip1(n21186), .ip2(n21136), .op(n21565) );
  nor3_1 U25229 ( .ip1(n21137), .ip2(n21577), .ip3(n21565), .op(n21184) );
  nor2_1 U25230 ( .ip1(\x[92][14] ), .ip2(n24327), .op(n21182) );
  and2_1 U25231 ( .ip1(n23895), .ip2(\x[92][13] ), .op(n21180) );
  inv_1 U25232 ( .ip(\x[92][12] ), .op(n21178) );
  nand2_1 U25233 ( .ip1(\x[92][11] ), .ip2(n24239), .op(n21140) );
  nand2_1 U25234 ( .ip1(\x[92][10] ), .ip2(n23146), .op(n21138) );
  nor2_1 U25235 ( .ip1(\x[92][11] ), .ip2(n24371), .op(n21169) );
  or2_1 U25236 ( .ip1(n21138), .ip2(n21169), .op(n21139) );
  nand2_1 U25237 ( .ip1(n21140), .ip2(n21139), .op(n21175) );
  inv_1 U25238 ( .ip(\x[92][9] ), .op(n21170) );
  nor2_1 U25239 ( .ip1(n21171), .ip2(n21170), .op(n21167) );
  inv_1 U25240 ( .ip(\x[92][7] ), .op(n21164) );
  nor2_1 U25241 ( .ip1(n17732), .ip2(n21164), .op(n21161) );
  inv_1 U25242 ( .ip(\x[92][5] ), .op(n21159) );
  inv_1 U25243 ( .ip(\x[92][4] ), .op(n21151) );
  nor2_1 U25244 ( .ip1(n24462), .ip2(n21151), .op(n21149) );
  inv_1 U25245 ( .ip(\x[92][3] ), .op(n21147) );
  inv_1 U25246 ( .ip(\x[92][1] ), .op(n21142) );
  nor2_1 U25247 ( .ip1(sig_in[1]), .ip2(n21142), .op(n21144) );
  inv_1 U25248 ( .ip(\x[92][0] ), .op(n21141) );
  not_ab_or_c_or_d U25249 ( .ip1(n24467), .ip2(n21142), .ip3(n23195), .ip4(
        n21141), .op(n21143) );
  not_ab_or_c_or_d U25250 ( .ip1(\x[92][2] ), .ip2(n24470), .ip3(n21144), 
        .ip4(n21143), .op(n21146) );
  nor2_1 U25251 ( .ip1(\x[92][2] ), .ip2(n23659), .op(n21145) );
  not_ab_or_c_or_d U25252 ( .ip1(sig_in[3]), .ip2(n21147), .ip3(n21146), .ip4(
        n21145), .op(n21148) );
  not_ab_or_c_or_d U25253 ( .ip1(\x[92][3] ), .ip2(n24476), .ip3(n21149), 
        .ip4(n21148), .op(n21150) );
  or2_1 U25254 ( .ip1(sig_in[4]), .ip2(n21150), .op(n21153) );
  or2_1 U25255 ( .ip1(n21151), .ip2(n21150), .op(n21152) );
  nand2_1 U25256 ( .ip1(n21153), .ip2(n21152), .op(n21154) );
  or2_1 U25257 ( .ip1(\x[92][5] ), .ip2(n21154), .op(n21156) );
  or2_1 U25258 ( .ip1(n24482), .ip2(n21154), .op(n21155) );
  nand2_1 U25259 ( .ip1(n21156), .ip2(n21155), .op(n21158) );
  nor2_1 U25260 ( .ip1(\x[92][6] ), .ip2(n23509), .op(n21157) );
  not_ab_or_c_or_d U25261 ( .ip1(sig_in[5]), .ip2(n21159), .ip3(n21158), .ip4(
        n21157), .op(n21160) );
  not_ab_or_c_or_d U25262 ( .ip1(\x[92][6] ), .ip2(n24045), .ip3(n21161), 
        .ip4(n21160), .op(n21163) );
  nor2_1 U25263 ( .ip1(\x[92][8] ), .ip2(n24491), .op(n21162) );
  not_ab_or_c_or_d U25264 ( .ip1(sig_in[7]), .ip2(n21164), .ip3(n21163), .ip4(
        n21162), .op(n21166) );
  and2_1 U25265 ( .ip1(n23804), .ip2(\x[92][8] ), .op(n21165) );
  nor3_1 U25266 ( .ip1(n21167), .ip2(n21166), .ip3(n21165), .op(n21173) );
  nor2_1 U25267 ( .ip1(\x[92][10] ), .ip2(n24457), .op(n21168) );
  ab_or_c_or_d U25268 ( .ip1(n21171), .ip2(n21170), .ip3(n21169), .ip4(n21168), 
        .op(n21172) );
  nor2_1 U25269 ( .ip1(n21173), .ip2(n21172), .op(n21174) );
  not_ab_or_c_or_d U25270 ( .ip1(\x[92][12] ), .ip2(n24449), .ip3(n21175), 
        .ip4(n21174), .op(n21177) );
  nor2_1 U25271 ( .ip1(\x[92][13] ), .ip2(n24376), .op(n21176) );
  not_ab_or_c_or_d U25272 ( .ip1(sig_in[12]), .ip2(n21178), .ip3(n21177), 
        .ip4(n21176), .op(n21179) );
  not_ab_or_c_or_d U25273 ( .ip1(\x[92][14] ), .ip2(n24382), .ip3(n21180), 
        .ip4(n21179), .op(n21181) );
  not_ab_or_c_or_d U25274 ( .ip1(\x[92][15] ), .ip2(n24180), .ip3(n21182), 
        .ip4(n21181), .op(n21557) );
  nor2_1 U25275 ( .ip1(\x[92][15] ), .ip2(n24180), .op(n21560) );
  nor2_1 U25276 ( .ip1(n21557), .ip2(n21560), .op(n21183) );
  not_ab_or_c_or_d U25277 ( .ip1(n21186), .ip2(n21185), .ip3(n21184), .ip4(
        n21183), .op(n24548) );
  nor2_1 U25278 ( .ip1(\x[94][15] ), .ip2(n24329), .op(n21266) );
  nand2_1 U25279 ( .ip1(n23143), .ip2(\x[94][15] ), .op(n21535) );
  inv_1 U25280 ( .ip(n21535), .op(n21190) );
  nor2_1 U25281 ( .ip1(\x[94][14] ), .ip2(n24327), .op(n21189) );
  nor2_1 U25282 ( .ip1(\x[94][13] ), .ip2(n24137), .op(n21188) );
  nor2_1 U25283 ( .ip1(\x[94][12] ), .ip2(n24079), .op(n21187) );
  nor4_1 U25284 ( .ip1(n21190), .ip2(n21189), .ip3(n21188), .ip4(n21187), .op(
        n21537) );
  nor2_1 U25285 ( .ip1(n21266), .ip2(n21537), .op(n21274) );
  nand2_1 U25286 ( .ip1(n24329), .ip2(\x[93][15] ), .op(n21232) );
  nand2_1 U25287 ( .ip1(n23938), .ip2(\x[93][14] ), .op(n21192) );
  or2_1 U25288 ( .ip1(n24384), .ip2(\x[93][15] ), .op(n21549) );
  nand2_1 U25289 ( .ip1(\x[93][13] ), .ip2(n24235), .op(n21191) );
  nand3_1 U25290 ( .ip1(n21192), .ip2(n21549), .ip3(n21191), .op(n21193) );
  inv_1 U25291 ( .ip(n21193), .op(n21559) );
  nand2_1 U25292 ( .ip1(\x[93][12] ), .ip2(n24233), .op(n21194) );
  nand2_1 U25293 ( .ip1(n21559), .ip2(n21194), .op(n21552) );
  and2_1 U25294 ( .ip1(n21232), .ip2(n21552), .op(n21273) );
  nor2_1 U25295 ( .ip1(\x[93][11] ), .ip2(n24371), .op(n21196) );
  nor2_1 U25296 ( .ip1(\x[93][10] ), .ip2(n24457), .op(n21195) );
  nor2_1 U25297 ( .ip1(n21196), .ip2(n21195), .op(n21228) );
  inv_1 U25298 ( .ip(n21228), .op(n21197) );
  nand2_1 U25299 ( .ip1(\x[93][11] ), .ip2(n24239), .op(n21202) );
  nand2_1 U25300 ( .ip1(n21197), .ip2(n21202), .op(n21554) );
  nand2_1 U25301 ( .ip1(\x[93][9] ), .ip2(n24164), .op(n21201) );
  nand2_1 U25302 ( .ip1(\x[93][10] ), .ip2(n23146), .op(n21200) );
  nor2_1 U25303 ( .ip1(n24455), .ip2(\x[93][9] ), .op(n21225) );
  inv_1 U25304 ( .ip(n21225), .op(n21198) );
  nand3_1 U25305 ( .ip1(\x[93][8] ), .ip2(n23971), .ip3(n21198), .op(n21199)
         );
  nand4_1 U25306 ( .ip1(n21202), .ip2(n21201), .ip3(n21200), .ip4(n21199), 
        .op(n21203) );
  nand2_1 U25307 ( .ip1(n21554), .ip2(n21203), .op(n21551) );
  not_ab_or_c_or_d U25308 ( .ip1(\x[93][7] ), .ip2(n24142), .ip3(\x[93][6] ), 
        .ip4(n23770), .op(n21227) );
  inv_1 U25309 ( .ip(\x[93][4] ), .op(n21217) );
  and2_1 U25310 ( .ip1(n23659), .ip2(\x[93][2] ), .op(n21209) );
  nand2_1 U25311 ( .ip1(\x[93][1] ), .ip2(n21685), .op(n21207) );
  nand2_1 U25312 ( .ip1(\x[93][0] ), .ip2(n24143), .op(n21206) );
  nor2_1 U25313 ( .ip1(\x[93][2] ), .ip2(n23717), .op(n21205) );
  nor2_1 U25314 ( .ip1(\x[93][1] ), .ip2(n20652), .op(n21204) );
  not_ab_or_c_or_d U25315 ( .ip1(n21207), .ip2(n21206), .ip3(n21205), .ip4(
        n21204), .op(n21208) );
  not_ab_or_c_or_d U25316 ( .ip1(\x[93][3] ), .ip2(n22525), .ip3(n21209), 
        .ip4(n21208), .op(n21211) );
  nor2_1 U25317 ( .ip1(\x[93][3] ), .ip2(n24342), .op(n21210) );
  nor2_1 U25318 ( .ip1(n21211), .ip2(n21210), .op(n21212) );
  or2_1 U25319 ( .ip1(\x[93][4] ), .ip2(n21212), .op(n21214) );
  or2_1 U25320 ( .ip1(n24347), .ip2(n21212), .op(n21213) );
  nand2_1 U25321 ( .ip1(n21214), .ip2(n21213), .op(n21216) );
  nor2_1 U25322 ( .ip1(\x[93][5] ), .ip2(n23283), .op(n21215) );
  not_ab_or_c_or_d U25323 ( .ip1(sig_in[4]), .ip2(n21217), .ip3(n21216), .ip4(
        n21215), .op(n21221) );
  nand2_1 U25324 ( .ip1(\x[93][7] ), .ip2(n24044), .op(n21219) );
  nand2_1 U25325 ( .ip1(\x[93][6] ), .ip2(n24485), .op(n21218) );
  nand2_1 U25326 ( .ip1(n21219), .ip2(n21218), .op(n21220) );
  not_ab_or_c_or_d U25327 ( .ip1(\x[93][5] ), .ip2(n24482), .ip3(n21221), 
        .ip4(n21220), .op(n21224) );
  nor2_1 U25328 ( .ip1(\x[93][8] ), .ip2(n24491), .op(n21223) );
  nor2_1 U25329 ( .ip1(\x[93][7] ), .ip2(n24044), .op(n21222) );
  or4_1 U25330 ( .ip1(n21225), .ip2(n21224), .ip3(n21223), .ip4(n21222), .op(
        n21226) );
  nor2_1 U25331 ( .ip1(n21227), .ip2(n21226), .op(n21555) );
  nand2_1 U25332 ( .ip1(n21228), .ip2(n21555), .op(n21233) );
  nor2_1 U25333 ( .ip1(\x[93][13] ), .ip2(n24137), .op(n21230) );
  nor2_1 U25334 ( .ip1(\x[93][12] ), .ip2(n24079), .op(n21229) );
  or2_1 U25335 ( .ip1(n21230), .ip2(n21229), .op(n21558) );
  or2_1 U25336 ( .ip1(n24185), .ip2(\x[93][14] ), .op(n21231) );
  nand2_1 U25337 ( .ip1(n21232), .ip2(n21231), .op(n21550) );
  not_ab_or_c_or_d U25338 ( .ip1(n21551), .ip2(n21233), .ip3(n21558), .ip4(
        n21550), .op(n21272) );
  and2_1 U25339 ( .ip1(n24451), .ip2(\x[94][10] ), .op(n21263) );
  inv_1 U25340 ( .ip(\x[94][9] ), .op(n21261) );
  inv_1 U25341 ( .ip(\x[94][8] ), .op(n21253) );
  nor2_1 U25342 ( .ip1(n21253), .ip2(sig_in[8]), .op(n21255) );
  and2_1 U25343 ( .ip1(n24461), .ip2(\x[94][7] ), .op(n21250) );
  inv_1 U25344 ( .ip(\x[94][3] ), .op(n21240) );
  nor2_1 U25345 ( .ip1(\x[94][2] ), .ip2(n23659), .op(n21239) );
  inv_1 U25346 ( .ip(\x[94][1] ), .op(n21235) );
  nor2_1 U25347 ( .ip1(n24464), .ip2(n21235), .op(n21237) );
  inv_1 U25348 ( .ip(\x[94][0] ), .op(n21234) );
  not_ab_or_c_or_d U25349 ( .ip1(n24467), .ip2(n21235), .ip3(n23195), .ip4(
        n21234), .op(n21236) );
  not_ab_or_c_or_d U25350 ( .ip1(\x[94][2] ), .ip2(n24470), .ip3(n21237), 
        .ip4(n21236), .op(n21238) );
  not_ab_or_c_or_d U25351 ( .ip1(sig_in[3]), .ip2(n21240), .ip3(n21239), .ip4(
        n21238), .op(n21244) );
  nand2_1 U25352 ( .ip1(\x[94][5] ), .ip2(n24119), .op(n21242) );
  nand2_1 U25353 ( .ip1(\x[94][4] ), .ip2(n23860), .op(n21241) );
  nand2_1 U25354 ( .ip1(n21242), .ip2(n21241), .op(n21243) );
  not_ab_or_c_or_d U25355 ( .ip1(\x[94][3] ), .ip2(n22525), .ip3(n21244), 
        .ip4(n21243), .op(n21248) );
  nor2_1 U25356 ( .ip1(\x[94][6] ), .ip2(n23770), .op(n21247) );
  nor2_1 U25357 ( .ip1(\x[94][5] ), .ip2(n23283), .op(n21246) );
  not_ab_or_c_or_d U25358 ( .ip1(\x[94][5] ), .ip2(n24482), .ip3(\x[94][4] ), 
        .ip4(n24256), .op(n21245) );
  nor4_1 U25359 ( .ip1(n21248), .ip2(n21247), .ip3(n21246), .ip4(n21245), .op(
        n21249) );
  not_ab_or_c_or_d U25360 ( .ip1(\x[94][6] ), .ip2(n24045), .ip3(n21250), 
        .ip4(n21249), .op(n21252) );
  nor2_1 U25361 ( .ip1(\x[94][7] ), .ip2(n24492), .op(n21251) );
  not_ab_or_c_or_d U25362 ( .ip1(sig_in[8]), .ip2(n21253), .ip3(n21252), .ip4(
        n21251), .op(n21254) );
  or2_1 U25363 ( .ip1(n21255), .ip2(n21254), .op(n21256) );
  or2_1 U25364 ( .ip1(\x[94][9] ), .ip2(n21256), .op(n21258) );
  or2_1 U25365 ( .ip1(n24269), .ip2(n21256), .op(n21257) );
  nand2_1 U25366 ( .ip1(n21258), .ip2(n21257), .op(n21260) );
  nor2_1 U25367 ( .ip1(\x[94][10] ), .ip2(n24457), .op(n21259) );
  not_ab_or_c_or_d U25368 ( .ip1(sig_in[9]), .ip2(n21261), .ip3(n21260), .ip4(
        n21259), .op(n21262) );
  not_ab_or_c_or_d U25369 ( .ip1(\x[94][11] ), .ip2(n24136), .ip3(n21263), 
        .ip4(n21262), .op(n21265) );
  nor2_1 U25370 ( .ip1(\x[94][11] ), .ip2(n24239), .op(n21264) );
  nor2_1 U25371 ( .ip1(n21265), .ip2(n21264), .op(n21536) );
  inv_1 U25372 ( .ip(n21266), .op(n21270) );
  nand2_1 U25373 ( .ip1(\x[94][12] ), .ip2(n24450), .op(n21269) );
  nand2_1 U25374 ( .ip1(\x[94][14] ), .ip2(n23938), .op(n21268) );
  nand2_1 U25375 ( .ip1(\x[94][13] ), .ip2(n24081), .op(n21267) );
  nand4_1 U25376 ( .ip1(n21270), .ip2(n21269), .ip3(n21268), .ip4(n21267), 
        .op(n21534) );
  nor2_1 U25377 ( .ip1(n21536), .ip2(n21534), .op(n21271) );
  nor4_1 U25378 ( .ip1(n21274), .ip2(n21273), .ip3(n21272), .ip4(n21271), .op(
        n24542) );
  nand2_1 U25379 ( .ip1(n24230), .ip2(\x[96][14] ), .op(n21277) );
  nor2_1 U25380 ( .ip1(n24384), .ip2(\x[96][15] ), .op(n21327) );
  inv_1 U25381 ( .ip(n21327), .op(n21276) );
  nand2_1 U25382 ( .ip1(\x[96][13] ), .ip2(n24235), .op(n21275) );
  nand3_1 U25383 ( .ip1(n21277), .ip2(n21276), .ip3(n21275), .op(n21323) );
  or2_1 U25384 ( .ip1(\x[96][12] ), .ip2(n21323), .op(n21279) );
  or2_1 U25385 ( .ip1(n24079), .ip2(n21323), .op(n21278) );
  nand2_1 U25386 ( .ip1(n21279), .ip2(n21278), .op(n21519) );
  nor2_1 U25387 ( .ip1(n24371), .ip2(\x[96][11] ), .op(n21317) );
  inv_1 U25388 ( .ip(\x[96][9] ), .op(n21313) );
  inv_1 U25389 ( .ip(\x[96][8] ), .op(n21305) );
  nor2_1 U25390 ( .ip1(n23779), .ip2(n21305), .op(n21303) );
  inv_1 U25391 ( .ip(\x[96][3] ), .op(n21286) );
  inv_1 U25392 ( .ip(\x[96][1] ), .op(n21281) );
  nor2_1 U25393 ( .ip1(n24464), .ip2(n21281), .op(n21283) );
  inv_1 U25394 ( .ip(\x[96][0] ), .op(n21280) );
  not_ab_or_c_or_d U25395 ( .ip1(n24467), .ip2(n21281), .ip3(n23195), .ip4(
        n21280), .op(n21282) );
  not_ab_or_c_or_d U25396 ( .ip1(\x[96][2] ), .ip2(n24107), .ip3(n21283), 
        .ip4(n21282), .op(n21285) );
  nor2_1 U25397 ( .ip1(\x[96][2] ), .ip2(n23659), .op(n21284) );
  not_ab_or_c_or_d U25398 ( .ip1(sig_in[3]), .ip2(n21286), .ip3(n21285), .ip4(
        n21284), .op(n21290) );
  nand2_1 U25399 ( .ip1(\x[96][5] ), .ip2(n24119), .op(n21288) );
  nand2_1 U25400 ( .ip1(\x[96][4] ), .ip2(n23721), .op(n21287) );
  nand2_1 U25401 ( .ip1(n21288), .ip2(n21287), .op(n21289) );
  not_ab_or_c_or_d U25402 ( .ip1(\x[96][3] ), .ip2(n24476), .ip3(n21290), 
        .ip4(n21289), .op(n21294) );
  nor2_1 U25403 ( .ip1(\x[96][5] ), .ip2(n23283), .op(n21293) );
  nor2_1 U25404 ( .ip1(\x[96][6] ), .ip2(n23770), .op(n21292) );
  not_ab_or_c_or_d U25405 ( .ip1(\x[96][5] ), .ip2(n24482), .ip3(\x[96][4] ), 
        .ip4(n24256), .op(n21291) );
  nor4_1 U25406 ( .ip1(n21294), .ip2(n21293), .ip3(n21292), .ip4(n21291), .op(
        n21295) );
  or2_1 U25407 ( .ip1(\x[96][6] ), .ip2(n21295), .op(n21297) );
  or2_1 U25408 ( .ip1(n24045), .ip2(n21295), .op(n21296) );
  nand2_1 U25409 ( .ip1(n21297), .ip2(n21296), .op(n21298) );
  or2_1 U25410 ( .ip1(sig_in[7]), .ip2(n21298), .op(n21301) );
  inv_1 U25411 ( .ip(\x[96][7] ), .op(n21299) );
  or2_1 U25412 ( .ip1(n21299), .ip2(n21298), .op(n21300) );
  nand2_1 U25413 ( .ip1(n21301), .ip2(n21300), .op(n21302) );
  not_ab_or_c_or_d U25414 ( .ip1(\x[96][7] ), .ip2(n24142), .ip3(n21303), 
        .ip4(n21302), .op(n21304) );
  or2_1 U25415 ( .ip1(n23779), .ip2(n21304), .op(n21307) );
  or2_1 U25416 ( .ip1(n21305), .ip2(n21304), .op(n21306) );
  nand2_1 U25417 ( .ip1(n21307), .ip2(n21306), .op(n21308) );
  or2_1 U25418 ( .ip1(\x[96][9] ), .ip2(n21308), .op(n21310) );
  or2_1 U25419 ( .ip1(n24269), .ip2(n21308), .op(n21309) );
  nand2_1 U25420 ( .ip1(n21310), .ip2(n21309), .op(n21312) );
  nor2_1 U25421 ( .ip1(\x[96][10] ), .ip2(n24457), .op(n21311) );
  not_ab_or_c_or_d U25422 ( .ip1(sig_in[9]), .ip2(n21313), .ip3(n21312), .ip4(
        n21311), .op(n21315) );
  and2_1 U25423 ( .ip1(n24451), .ip2(\x[96][10] ), .op(n21314) );
  not_ab_or_c_or_d U25424 ( .ip1(\x[96][11] ), .ip2(n24136), .ip3(n21315), 
        .ip4(n21314), .op(n21316) );
  nor2_1 U25425 ( .ip1(n21317), .ip2(n21316), .op(n21529) );
  inv_1 U25426 ( .ip(n21529), .op(n21373) );
  and2_1 U25427 ( .ip1(n23895), .ip2(\x[95][13] ), .op(n21318) );
  nor2_1 U25428 ( .ip1(\x[95][15] ), .ip2(n24180), .op(n21533) );
  not_ab_or_c_or_d U25429 ( .ip1(\x[95][14] ), .ip2(n24382), .ip3(n21318), 
        .ip4(n21533), .op(n21543) );
  and2_1 U25430 ( .ip1(n24186), .ip2(\x[95][15] ), .op(n21364) );
  or2_1 U25431 ( .ip1(n21543), .ip2(n21364), .op(n21320) );
  nand2_1 U25432 ( .ip1(\x[95][12] ), .ip2(n24450), .op(n21539) );
  or2_1 U25433 ( .ip1(n21539), .ip2(n21364), .op(n21319) );
  nand2_1 U25434 ( .ip1(n21320), .ip2(n21319), .op(n21372) );
  nor2_1 U25435 ( .ip1(\x[96][13] ), .ip2(n24376), .op(n21322) );
  nor2_1 U25436 ( .ip1(\x[96][12] ), .ip2(n24079), .op(n21321) );
  nor2_1 U25437 ( .ip1(n21322), .ip2(n21321), .op(n21528) );
  or2_1 U25438 ( .ip1(n21528), .ip2(n21323), .op(n21370) );
  nor2_1 U25439 ( .ip1(\x[96][14] ), .ip2(n24327), .op(n21324) );
  or2_1 U25440 ( .ip1(\x[96][15] ), .ip2(n21324), .op(n21326) );
  or2_1 U25441 ( .ip1(n24384), .ip2(n21324), .op(n21325) );
  nand2_1 U25442 ( .ip1(n21326), .ip2(n21325), .op(n21527) );
  nor2_1 U25443 ( .ip1(n21527), .ip2(n21327), .op(n21518) );
  inv_1 U25444 ( .ip(n21518), .op(n21369) );
  inv_1 U25445 ( .ip(\x[95][10] ), .op(n21352) );
  nor2_1 U25446 ( .ip1(n21352), .ip2(sig_in[10]), .op(n21354) );
  nor2_1 U25447 ( .ip1(\x[95][9] ), .ip2(n24164), .op(n21351) );
  and2_1 U25448 ( .ip1(n23804), .ip2(\x[95][8] ), .op(n21349) );
  inv_1 U25449 ( .ip(\x[95][7] ), .op(n21347) );
  nor2_1 U25450 ( .ip1(sig_in[7]), .ip2(n21347), .op(n21344) );
  inv_1 U25451 ( .ip(\x[95][3] ), .op(n21334) );
  inv_1 U25452 ( .ip(\x[95][1] ), .op(n21329) );
  nor2_1 U25453 ( .ip1(n24464), .ip2(n21329), .op(n21331) );
  inv_1 U25454 ( .ip(\x[95][0] ), .op(n21328) );
  not_ab_or_c_or_d U25455 ( .ip1(n22513), .ip2(n21329), .ip3(n23195), .ip4(
        n21328), .op(n21330) );
  not_ab_or_c_or_d U25456 ( .ip1(\x[95][2] ), .ip2(n24470), .ip3(n21331), 
        .ip4(n21330), .op(n21333) );
  nor2_1 U25457 ( .ip1(\x[95][2] ), .ip2(n23659), .op(n21332) );
  not_ab_or_c_or_d U25458 ( .ip1(sig_in[3]), .ip2(n21334), .ip3(n21333), .ip4(
        n21332), .op(n21338) );
  nand2_1 U25459 ( .ip1(\x[95][5] ), .ip2(n24119), .op(n21336) );
  nand2_1 U25460 ( .ip1(\x[95][4] ), .ip2(n23721), .op(n21335) );
  nand2_1 U25461 ( .ip1(n21336), .ip2(n21335), .op(n21337) );
  not_ab_or_c_or_d U25462 ( .ip1(\x[95][3] ), .ip2(n22525), .ip3(n21338), 
        .ip4(n21337), .op(n21342) );
  nor2_1 U25463 ( .ip1(\x[95][6] ), .ip2(n23509), .op(n21341) );
  nor2_1 U25464 ( .ip1(\x[95][5] ), .ip2(n23283), .op(n21340) );
  not_ab_or_c_or_d U25465 ( .ip1(\x[95][5] ), .ip2(n23600), .ip3(\x[95][4] ), 
        .ip4(n24347), .op(n21339) );
  nor4_1 U25466 ( .ip1(n21342), .ip2(n21341), .ip3(n21340), .ip4(n21339), .op(
        n21343) );
  not_ab_or_c_or_d U25467 ( .ip1(\x[95][6] ), .ip2(n24045), .ip3(n21344), 
        .ip4(n21343), .op(n21346) );
  nor2_1 U25468 ( .ip1(\x[95][8] ), .ip2(n24358), .op(n21345) );
  not_ab_or_c_or_d U25469 ( .ip1(sig_in[7]), .ip2(n21347), .ip3(n21346), .ip4(
        n21345), .op(n21348) );
  not_ab_or_c_or_d U25470 ( .ip1(\x[95][9] ), .ip2(n23981), .ip3(n21349), 
        .ip4(n21348), .op(n21350) );
  not_ab_or_c_or_d U25471 ( .ip1(sig_in[10]), .ip2(n21352), .ip3(n21351), 
        .ip4(n21350), .op(n21353) );
  or2_1 U25472 ( .ip1(n21354), .ip2(n21353), .op(n21355) );
  or2_1 U25473 ( .ip1(\x[95][11] ), .ip2(n21355), .op(n21357) );
  or2_1 U25474 ( .ip1(n24136), .ip2(n21355), .op(n21356) );
  nand2_1 U25475 ( .ip1(n21357), .ip2(n21356), .op(n21359) );
  nor2_1 U25476 ( .ip1(\x[95][11] ), .ip2(n24371), .op(n21358) );
  nor2_1 U25477 ( .ip1(n21359), .ip2(n21358), .op(n21538) );
  nor2_1 U25478 ( .ip1(\x[95][13] ), .ip2(n24332), .op(n21360) );
  or2_1 U25479 ( .ip1(sig_in[12]), .ip2(n21360), .op(n21363) );
  inv_1 U25480 ( .ip(\x[95][12] ), .op(n21361) );
  or2_1 U25481 ( .ip1(n21361), .ip2(n21360), .op(n21362) );
  nand2_1 U25482 ( .ip1(n21363), .ip2(n21362), .op(n21541) );
  or2_1 U25483 ( .ip1(sig_in[14]), .ip2(n21364), .op(n21367) );
  inv_1 U25484 ( .ip(\x[95][14] ), .op(n21365) );
  or2_1 U25485 ( .ip1(n21365), .ip2(n21364), .op(n21366) );
  nand2_1 U25486 ( .ip1(n21367), .ip2(n21366), .op(n21532) );
  nand3_1 U25487 ( .ip1(n21538), .ip2(n21541), .ip3(n21532), .op(n21368) );
  nand3_1 U25488 ( .ip1(n21370), .ip2(n21369), .ip3(n21368), .op(n21371) );
  not_ab_or_c_or_d U25489 ( .ip1(n21519), .ip2(n21373), .ip3(n21372), .ip4(
        n21371), .op(n24532) );
  nand2_1 U25490 ( .ip1(\x[97][15] ), .ip2(n24186), .op(n21465) );
  and2_1 U25491 ( .ip1(n23895), .ip2(\x[97][13] ), .op(n21374) );
  nor2_1 U25492 ( .ip1(\x[97][15] ), .ip2(n24180), .op(n21521) );
  not_ab_or_c_or_d U25493 ( .ip1(\x[97][14] ), .ip2(n24382), .ip3(n21374), 
        .ip4(n21521), .op(n21526) );
  nand2_1 U25494 ( .ip1(\x[97][12] ), .ip2(n24450), .op(n21514) );
  nand2_1 U25495 ( .ip1(n21526), .ip2(n21514), .op(n21464) );
  and2_1 U25496 ( .ip1(n24451), .ip2(\x[97][10] ), .op(n21399) );
  nor2_1 U25497 ( .ip1(\x[97][7] ), .ip2(n24044), .op(n21389) );
  inv_1 U25498 ( .ip(\x[97][6] ), .op(n21375) );
  nor3_1 U25499 ( .ip1(sig_in[6]), .ip2(n21389), .ip3(n21375), .op(n21392) );
  and2_1 U25500 ( .ip1(n24119), .ip2(\x[97][5] ), .op(n21386) );
  inv_1 U25501 ( .ip(\x[97][3] ), .op(n21384) );
  and2_1 U25502 ( .ip1(n24107), .ip2(\x[97][2] ), .op(n21381) );
  nand2_1 U25503 ( .ip1(\x[97][1] ), .ip2(n21685), .op(n21379) );
  nand2_1 U25504 ( .ip1(\x[97][0] ), .ip2(n24143), .op(n21378) );
  nor2_1 U25505 ( .ip1(\x[97][2] ), .ip2(n23717), .op(n21377) );
  nor2_1 U25506 ( .ip1(\x[97][1] ), .ip2(n21685), .op(n21376) );
  not_ab_or_c_or_d U25507 ( .ip1(n21379), .ip2(n21378), .ip3(n21377), .ip4(
        n21376), .op(n21380) );
  not_ab_or_c_or_d U25508 ( .ip1(\x[97][3] ), .ip2(n22525), .ip3(n21381), 
        .ip4(n21380), .op(n21383) );
  nor2_1 U25509 ( .ip1(\x[97][4] ), .ip2(n24347), .op(n21382) );
  not_ab_or_c_or_d U25510 ( .ip1(sig_in[3]), .ip2(n21384), .ip3(n21383), .ip4(
        n21382), .op(n21385) );
  not_ab_or_c_or_d U25511 ( .ip1(\x[97][4] ), .ip2(n23860), .ip3(n21386), 
        .ip4(n21385), .op(n21390) );
  nor2_1 U25512 ( .ip1(\x[97][6] ), .ip2(n23509), .op(n21388) );
  nor2_1 U25513 ( .ip1(\x[97][5] ), .ip2(n23283), .op(n21387) );
  nor4_1 U25514 ( .ip1(n21390), .ip2(n21389), .ip3(n21388), .ip4(n21387), .op(
        n21391) );
  not_ab_or_c_or_d U25515 ( .ip1(\x[97][8] ), .ip2(n24100), .ip3(n21392), 
        .ip4(n21391), .op(n21396) );
  nand2_1 U25516 ( .ip1(\x[97][7] ), .ip2(n24492), .op(n21395) );
  nor2_1 U25517 ( .ip1(\x[97][8] ), .ip2(n24358), .op(n21394) );
  nor2_1 U25518 ( .ip1(\x[97][9] ), .ip2(n24455), .op(n21393) );
  not_ab_or_c_or_d U25519 ( .ip1(n21396), .ip2(n21395), .ip3(n21394), .ip4(
        n21393), .op(n21398) );
  and2_1 U25520 ( .ip1(n23981), .ip2(\x[97][9] ), .op(n21397) );
  nor3_1 U25521 ( .ip1(n21399), .ip2(n21398), .ip3(n21397), .op(n21403) );
  nor2_1 U25522 ( .ip1(\x[97][11] ), .ip2(n24371), .op(n21401) );
  nor2_1 U25523 ( .ip1(\x[97][10] ), .ip2(n24457), .op(n21400) );
  or2_1 U25524 ( .ip1(n21401), .ip2(n21400), .op(n21402) );
  nor2_1 U25525 ( .ip1(n21403), .ip2(n21402), .op(n21404) );
  or2_1 U25526 ( .ip1(\x[97][11] ), .ip2(n21404), .op(n21406) );
  or2_1 U25527 ( .ip1(n24136), .ip2(n21404), .op(n21405) );
  nand2_1 U25528 ( .ip1(n21406), .ip2(n21405), .op(n21515) );
  or2_1 U25529 ( .ip1(n24185), .ip2(\x[97][14] ), .op(n21407) );
  nand2_1 U25530 ( .ip1(n21407), .ip2(n21465), .op(n21520) );
  nor2_1 U25531 ( .ip1(\x[97][13] ), .ip2(n24137), .op(n21409) );
  nor2_1 U25532 ( .ip1(\x[97][12] ), .ip2(n24449), .op(n21408) );
  nor2_1 U25533 ( .ip1(n21409), .ip2(n21408), .op(n21517) );
  inv_1 U25534 ( .ip(n21517), .op(n21410) );
  nor3_1 U25535 ( .ip1(n21515), .ip2(n21520), .ip3(n21410), .op(n21463) );
  and2_1 U25536 ( .ip1(n24332), .ip2(\x[98][13] ), .op(n21411) );
  nor2_1 U25537 ( .ip1(\x[98][15] ), .ip2(n24180), .op(n21457) );
  not_ab_or_c_or_d U25538 ( .ip1(\x[98][14] ), .ip2(n24382), .ip3(n21411), 
        .ip4(n21457), .op(n21461) );
  nor2_1 U25539 ( .ip1(\x[98][13] ), .ip2(n24376), .op(n21413) );
  nor2_1 U25540 ( .ip1(\x[98][12] ), .ip2(n24449), .op(n21412) );
  nor2_1 U25541 ( .ip1(n21413), .ip2(n21412), .op(n21467) );
  inv_1 U25542 ( .ip(n21467), .op(n21460) );
  nand2_1 U25543 ( .ip1(\x[98][10] ), .ip2(n23146), .op(n21443) );
  nor2_1 U25544 ( .ip1(\x[98][9] ), .ip2(n24164), .op(n21438) );
  inv_1 U25545 ( .ip(\x[98][8] ), .op(n21414) );
  nor3_1 U25546 ( .ip1(sig_in[8]), .ip2(n21438), .ip3(n21414), .op(n21441) );
  and2_1 U25547 ( .ip1(n24461), .ip2(\x[98][7] ), .op(n21435) );
  and2_1 U25548 ( .ip1(n24350), .ip2(\x[98][5] ), .op(n21415) );
  or2_1 U25549 ( .ip1(\x[98][4] ), .ip2(n21415), .op(n21417) );
  or2_1 U25550 ( .ip1(n23860), .ip2(n21415), .op(n21416) );
  nand2_1 U25551 ( .ip1(n21417), .ip2(n21416), .op(n21433) );
  nand2_1 U25552 ( .ip1(\x[98][1] ), .ip2(n21685), .op(n21420) );
  or2_1 U25553 ( .ip1(\x[98][1] ), .ip2(n21685), .op(n21418) );
  nand3_1 U25554 ( .ip1(n24143), .ip2(\x[98][0] ), .ip3(n21418), .op(n21419)
         );
  nand2_1 U25555 ( .ip1(n21420), .ip2(n21419), .op(n21421) );
  or2_1 U25556 ( .ip1(\x[98][2] ), .ip2(n21421), .op(n21423) );
  or2_1 U25557 ( .ip1(n24470), .ip2(n21421), .op(n21422) );
  nand2_1 U25558 ( .ip1(n21423), .ip2(n21422), .op(n21425) );
  nor2_1 U25559 ( .ip1(\x[98][2] ), .ip2(n23659), .op(n21424) );
  nor2_1 U25560 ( .ip1(n21425), .ip2(n21424), .op(n21426) );
  nand2_1 U25561 ( .ip1(n21426), .ip2(\x[98][3] ), .op(n21429) );
  nor2_1 U25562 ( .ip1(\x[98][4] ), .ip2(n23721), .op(n21428) );
  nor2_1 U25563 ( .ip1(n21426), .ip2(\x[98][3] ), .op(n21427) );
  ab_or_c_or_d U25564 ( .ip1(sig_in[3]), .ip2(n21429), .ip3(n21428), .ip4(
        n21427), .op(n21432) );
  nor2_1 U25565 ( .ip1(\x[98][6] ), .ip2(n23509), .op(n21431) );
  nor2_1 U25566 ( .ip1(\x[98][5] ), .ip2(n23283), .op(n21430) );
  not_ab_or_c_or_d U25567 ( .ip1(n21433), .ip2(n21432), .ip3(n21431), .ip4(
        n21430), .op(n21434) );
  not_ab_or_c_or_d U25568 ( .ip1(\x[98][6] ), .ip2(n23770), .ip3(n21435), 
        .ip4(n21434), .op(n21439) );
  nor2_1 U25569 ( .ip1(\x[98][8] ), .ip2(n24358), .op(n21437) );
  nor2_1 U25570 ( .ip1(\x[98][7] ), .ip2(n24492), .op(n21436) );
  nor4_1 U25571 ( .ip1(n21439), .ip2(n21438), .ip3(n21437), .ip4(n21436), .op(
        n21440) );
  not_ab_or_c_or_d U25572 ( .ip1(\x[98][9] ), .ip2(n23981), .ip3(n21441), 
        .ip4(n21440), .op(n21442) );
  nand2_1 U25573 ( .ip1(n21443), .ip2(n21442), .op(n21449) );
  nor2_1 U25574 ( .ip1(\x[98][10] ), .ip2(n24457), .op(n21444) );
  or2_1 U25575 ( .ip1(sig_in[11]), .ip2(n21444), .op(n21447) );
  inv_1 U25576 ( .ip(\x[98][11] ), .op(n21445) );
  or2_1 U25577 ( .ip1(n21445), .ip2(n21444), .op(n21446) );
  nand2_1 U25578 ( .ip1(n21447), .ip2(n21446), .op(n21448) );
  nand2_1 U25579 ( .ip1(n21449), .ip2(n21448), .op(n21451) );
  nand2_1 U25580 ( .ip1(\x[98][11] ), .ip2(n21793), .op(n21450) );
  nand2_1 U25581 ( .ip1(n21451), .ip2(n21450), .op(n21468) );
  nand2_1 U25582 ( .ip1(\x[98][12] ), .ip2(n24450), .op(n21452) );
  nand2_1 U25583 ( .ip1(n21461), .ip2(n21452), .op(n21513) );
  nor2_1 U25584 ( .ip1(n21468), .ip2(n21513), .op(n21459) );
  nand2_1 U25585 ( .ip1(n23143), .ip2(\x[98][15] ), .op(n21512) );
  inv_1 U25586 ( .ip(n21512), .op(n21453) );
  or2_1 U25587 ( .ip1(sig_in[14]), .ip2(n21453), .op(n21456) );
  inv_1 U25588 ( .ip(\x[98][14] ), .op(n21454) );
  or2_1 U25589 ( .ip1(n21454), .ip2(n21453), .op(n21455) );
  nand2_1 U25590 ( .ip1(n21456), .ip2(n21455), .op(n21466) );
  nor2_1 U25591 ( .ip1(n21457), .ip2(n21466), .op(n21458) );
  ab_or_c_or_d U25592 ( .ip1(n21461), .ip2(n21460), .ip3(n21459), .ip4(n21458), 
        .op(n21462) );
  not_ab_or_c_or_d U25593 ( .ip1(n21465), .ip2(n21464), .ip3(n21463), .ip4(
        n21462), .op(n27336) );
  and3_1 U25594 ( .ip1(n21468), .ip2(n21467), .ip3(n21466), .op(n21511) );
  nand2_1 U25595 ( .ip1(\x[99][11] ), .ip2(n24239), .op(n21471) );
  nand2_1 U25596 ( .ip1(\x[99][10] ), .ip2(n23146), .op(n21469) );
  nor2_1 U25597 ( .ip1(\x[99][11] ), .ip2(n24371), .op(n21472) );
  or2_1 U25598 ( .ip1(n21469), .ip2(n21472), .op(n21470) );
  nand2_1 U25599 ( .ip1(n21471), .ip2(n21470), .op(n21503) );
  nand2_1 U25600 ( .ip1(n24449), .ip2(\x[99][12] ), .op(n21501) );
  or2_1 U25601 ( .ip1(n20880), .ip2(\x[99][10] ), .op(n21498) );
  inv_1 U25602 ( .ip(\x[99][9] ), .op(n21474) );
  not_ab_or_c_or_d U25603 ( .ip1(\x[99][9] ), .ip2(n24164), .ip3(\x[99][8] ), 
        .ip4(n24358), .op(n21473) );
  not_ab_or_c_or_d U25604 ( .ip1(sig_in[9]), .ip2(n21474), .ip3(n21473), .ip4(
        n21472), .op(n21497) );
  nand2_1 U25605 ( .ip1(\x[99][8] ), .ip2(n24491), .op(n21495) );
  nand2_1 U25606 ( .ip1(\x[99][7] ), .ip2(n24492), .op(n21494) );
  nand2_1 U25607 ( .ip1(\x[99][9] ), .ip2(n24269), .op(n21493) );
  and2_1 U25608 ( .ip1(n23283), .ip2(\x[99][5] ), .op(n21483) );
  inv_1 U25609 ( .ip(\x[99][3] ), .op(n21481) );
  nor2_1 U25610 ( .ip1(\x[99][2] ), .ip2(n23659), .op(n21480) );
  inv_1 U25611 ( .ip(\x[99][1] ), .op(n21476) );
  nor2_1 U25612 ( .ip1(sig_in[1]), .ip2(n21476), .op(n21478) );
  inv_1 U25613 ( .ip(\x[99][0] ), .op(n21475) );
  not_ab_or_c_or_d U25614 ( .ip1(n22513), .ip2(n21476), .ip3(n23195), .ip4(
        n21475), .op(n21477) );
  not_ab_or_c_or_d U25615 ( .ip1(\x[99][2] ), .ip2(n24107), .ip3(n21478), 
        .ip4(n21477), .op(n21479) );
  not_ab_or_c_or_d U25616 ( .ip1(sig_in[3]), .ip2(n21481), .ip3(n21480), .ip4(
        n21479), .op(n21482) );
  not_ab_or_c_or_d U25617 ( .ip1(\x[99][3] ), .ip2(n24476), .ip3(n21483), 
        .ip4(n21482), .op(n21487) );
  nand2_1 U25618 ( .ip1(\x[99][4] ), .ip2(n24347), .op(n21486) );
  not_ab_or_c_or_d U25619 ( .ip1(\x[99][5] ), .ip2(n24482), .ip3(\x[99][4] ), 
        .ip4(n24256), .op(n21485) );
  nor2_1 U25620 ( .ip1(\x[99][5] ), .ip2(n23283), .op(n21484) );
  not_ab_or_c_or_d U25621 ( .ip1(n21487), .ip2(n21486), .ip3(n21485), .ip4(
        n21484), .op(n21488) );
  nand2_1 U25622 ( .ip1(n21488), .ip2(\x[99][6] ), .op(n21491) );
  nor2_1 U25623 ( .ip1(\x[99][7] ), .ip2(n24044), .op(n21490) );
  nor2_1 U25624 ( .ip1(n21488), .ip2(\x[99][6] ), .op(n21489) );
  ab_or_c_or_d U25625 ( .ip1(sig_in[6]), .ip2(n21491), .ip3(n21490), .ip4(
        n21489), .op(n21492) );
  nand4_1 U25626 ( .ip1(n21495), .ip2(n21494), .ip3(n21493), .ip4(n21492), 
        .op(n21496) );
  nand3_1 U25627 ( .ip1(n21498), .ip2(n21497), .ip3(n21496), .op(n21500) );
  nand2_1 U25628 ( .ip1(\x[99][13] ), .ip2(n24235), .op(n21499) );
  nand3_1 U25629 ( .ip1(n21501), .ip2(n21500), .ip3(n21499), .op(n21502) );
  not_ab_or_c_or_d U25630 ( .ip1(\x[99][14] ), .ip2(n24382), .ip3(n21503), 
        .ip4(n21502), .op(n21508) );
  inv_1 U25631 ( .ip(\x[99][14] ), .op(n21506) );
  nor2_1 U25632 ( .ip1(\x[99][13] ), .ip2(n24376), .op(n21505) );
  nor2_1 U25633 ( .ip1(\x[99][12] ), .ip2(n24450), .op(n21504) );
  ab_or_c_or_d U25634 ( .ip1(sig_in[14]), .ip2(n21506), .ip3(n21505), .ip4(
        n21504), .op(n21507) );
  not_ab_or_c_or_d U25635 ( .ip1(\x[99][15] ), .ip2(n24384), .ip3(n21508), 
        .ip4(n21507), .op(n21510) );
  nor2_1 U25636 ( .ip1(\x[99][15] ), .ip2(n24329), .op(n21509) );
  nor2_1 U25637 ( .ip1(n21510), .ip2(n21509), .op(n22385) );
  not_ab_or_c_or_d U25638 ( .ip1(n21513), .ip2(n21512), .ip3(n21511), .ip4(
        n22385), .op(n27335) );
  nor2_1 U25639 ( .ip1(n27336), .ip2(n27335), .op(n24529) );
  nand2_1 U25640 ( .ip1(n21515), .ip2(n21514), .op(n21516) );
  nand2_1 U25641 ( .ip1(n21517), .ip2(n21516), .op(n21525) );
  nor2_1 U25642 ( .ip1(n21519), .ip2(n21518), .op(n21524) );
  inv_1 U25643 ( .ip(n21520), .op(n21522) );
  nor2_1 U25644 ( .ip1(n21522), .ip2(n21521), .op(n21523) );
  not_ab_or_c_or_d U25645 ( .ip1(n21526), .ip2(n21525), .ip3(n21524), .ip4(
        n21523), .op(n21531) );
  nand3_1 U25646 ( .ip1(n21529), .ip2(n21528), .ip3(n21527), .op(n21530) );
  nand2_1 U25647 ( .ip1(n21531), .ip2(n21530), .op(n24530) );
  nand2_1 U25648 ( .ip1(n24529), .ip2(n24530), .op(n24534) );
  nor2_1 U25649 ( .ip1(n24532), .ip2(n24534), .op(n24535) );
  or2_1 U25650 ( .ip1(n21533), .ip2(n21532), .op(n21548) );
  nand2_1 U25651 ( .ip1(n21535), .ip2(n21534), .op(n21547) );
  nand2_1 U25652 ( .ip1(n21537), .ip2(n21536), .op(n21546) );
  inv_1 U25653 ( .ip(n21538), .op(n21540) );
  nand2_1 U25654 ( .ip1(n21540), .ip2(n21539), .op(n21542) );
  nand2_1 U25655 ( .ip1(n21542), .ip2(n21541), .op(n21544) );
  nand2_1 U25656 ( .ip1(n21544), .ip2(n21543), .op(n21545) );
  nand4_1 U25657 ( .ip1(n21548), .ip2(n21547), .ip3(n21546), .ip4(n21545), 
        .op(n24536) );
  nand2_1 U25658 ( .ip1(n24535), .ip2(n24536), .op(n24544) );
  nor2_1 U25659 ( .ip1(n24542), .ip2(n24544), .op(n24545) );
  nand2_1 U25660 ( .ip1(n21550), .ip2(n21549), .op(n21563) );
  inv_1 U25661 ( .ip(n21551), .op(n21553) );
  not_ab_or_c_or_d U25662 ( .ip1(n21555), .ip2(n21554), .ip3(n21553), .ip4(
        n21552), .op(n21556) );
  not_ab_or_c_or_d U25663 ( .ip1(n21559), .ip2(n21558), .ip3(n21557), .ip4(
        n21556), .op(n21562) );
  inv_1 U25664 ( .ip(n21560), .op(n21561) );
  nand3_1 U25665 ( .ip1(n21563), .ip2(n21562), .ip3(n21561), .op(n24546) );
  nand2_1 U25666 ( .ip1(n24545), .ip2(n24546), .op(n24549) );
  nor2_1 U25667 ( .ip1(n24548), .ip2(n24549), .op(n24559) );
  inv_1 U25668 ( .ip(n21564), .op(n21566) );
  nand2_1 U25669 ( .ip1(n21566), .ip2(n21565), .op(n21589) );
  or2_1 U25670 ( .ip1(n21568), .ip2(n21567), .op(n21588) );
  nor2_1 U25671 ( .ip1(n21570), .ip2(n21569), .op(n21571) );
  not_ab_or_c_or_d U25672 ( .ip1(n21574), .ip2(n21573), .ip3(n21572), .ip4(
        n21571), .op(n21576) );
  nand2_1 U25673 ( .ip1(n21576), .ip2(n21575), .op(n21581) );
  or2_1 U25674 ( .ip1(n21578), .ip2(n21577), .op(n21580) );
  nand3_1 U25675 ( .ip1(n21581), .ip2(n21580), .ip3(n21579), .op(n21587) );
  inv_1 U25676 ( .ip(n21582), .op(n21583) );
  nand3_1 U25677 ( .ip1(n21585), .ip2(n21584), .ip3(n21583), .op(n21586) );
  nand4_1 U25678 ( .ip1(n21589), .ip2(n21588), .ip3(n21587), .ip4(n21586), 
        .op(n24561) );
  nand2_1 U25679 ( .ip1(n24559), .ip2(n24561), .op(n24558) );
  nor2_1 U25680 ( .ip1(n24556), .ip2(n24558), .op(n24562) );
  not_ab_or_c_or_d U25681 ( .ip1(n21593), .ip2(n21592), .ip3(n21591), .ip4(
        n21590), .op(n21609) );
  inv_1 U25682 ( .ip(n21594), .op(n21595) );
  nand3_1 U25683 ( .ip1(n21597), .ip2(n21596), .ip3(n21595), .op(n21608) );
  inv_1 U25684 ( .ip(n21598), .op(n21599) );
  nand2_1 U25685 ( .ip1(n21600), .ip2(n21599), .op(n21607) );
  inv_1 U25686 ( .ip(n21601), .op(n21603) );
  nand2_1 U25687 ( .ip1(n21603), .ip2(n21602), .op(n21604) );
  nand2_1 U25688 ( .ip1(n21605), .ip2(n21604), .op(n21606) );
  nand4_1 U25689 ( .ip1(n21609), .ip2(n21608), .ip3(n21607), .ip4(n21606), 
        .op(n24563) );
  nand2_1 U25690 ( .ip1(n24562), .ip2(n24563), .op(n24528) );
  nor2_1 U25691 ( .ip1(n24526), .ip2(n24528), .op(n24572) );
  inv_1 U25692 ( .ip(n21610), .op(n21611) );
  nor2_1 U25693 ( .ip1(n21612), .ip2(n21611), .op(n21613) );
  not_ab_or_c_or_d U25694 ( .ip1(n21616), .ip2(n21615), .ip3(n21614), .ip4(
        n21613), .op(n21627) );
  nand3_1 U25695 ( .ip1(n21618), .ip2(n21617), .ip3(n21616), .op(n21626) );
  or2_1 U25696 ( .ip1(n21620), .ip2(n21619), .op(n21625) );
  inv_1 U25697 ( .ip(n21621), .op(n21622) );
  nand2_1 U25698 ( .ip1(n21623), .ip2(n21622), .op(n21624) );
  nand4_1 U25699 ( .ip1(n21627), .ip2(n21626), .ip3(n21625), .ip4(n21624), 
        .op(n24573) );
  nand2_1 U25700 ( .ip1(n24572), .ip2(n24573), .op(n24571) );
  and2_1 U25701 ( .ip1(n23895), .ip2(\x[101][13] ), .op(n21628) );
  nor2_1 U25702 ( .ip1(\x[101][15] ), .ip2(n24180), .op(n21640) );
  not_ab_or_c_or_d U25703 ( .ip1(\x[101][14] ), .ip2(n24382), .ip3(n21628), 
        .ip4(n21640), .op(n21717) );
  nor2_1 U25704 ( .ip1(\x[101][13] ), .ip2(n24376), .op(n21630) );
  nor2_1 U25705 ( .ip1(\x[101][12] ), .ip2(n24233), .op(n21629) );
  nor2_1 U25706 ( .ip1(n21630), .ip2(n21629), .op(n22378) );
  inv_1 U25707 ( .ip(n22378), .op(n21716) );
  and2_1 U25708 ( .ip1(n24332), .ip2(\x[100][13] ), .op(n21631) );
  or2_1 U25709 ( .ip1(\x[100][12] ), .ip2(n21631), .op(n21633) );
  or2_1 U25710 ( .ip1(n24079), .ip2(n21631), .op(n21632) );
  nand2_1 U25711 ( .ip1(n21633), .ip2(n21632), .op(n22387) );
  nand2_1 U25712 ( .ip1(n24329), .ip2(\x[100][15] ), .op(n21708) );
  inv_1 U25713 ( .ip(n21708), .op(n21634) );
  or2_1 U25714 ( .ip1(n22387), .ip2(n21634), .op(n21636) );
  nand2_1 U25715 ( .ip1(\x[100][14] ), .ip2(n24327), .op(n22394) );
  or2_1 U25716 ( .ip1(n22394), .ip2(n21634), .op(n21635) );
  nand2_1 U25717 ( .ip1(n21636), .ip2(n21635), .op(n21715) );
  nor2_1 U25718 ( .ip1(\x[101][14] ), .ip2(n24327), .op(n21637) );
  or2_1 U25719 ( .ip1(\x[101][15] ), .ip2(n21637), .op(n21639) );
  or2_1 U25720 ( .ip1(n24329), .ip2(n21637), .op(n21638) );
  nand2_1 U25721 ( .ip1(n21639), .ip2(n21638), .op(n22380) );
  nor2_1 U25722 ( .ip1(n21640), .ip2(n22380), .op(n22367) );
  nand2_1 U25723 ( .ip1(\x[101][9] ), .ip2(n24164), .op(n21666) );
  nor2_1 U25724 ( .ip1(\x[101][9] ), .ip2(n23981), .op(n21661) );
  inv_1 U25725 ( .ip(\x[101][8] ), .op(n21641) );
  nor3_1 U25726 ( .ip1(sig_in[8]), .ip2(n21661), .ip3(n21641), .op(n21664) );
  and2_1 U25727 ( .ip1(n24461), .ip2(\x[101][7] ), .op(n21658) );
  inv_1 U25728 ( .ip(\x[101][3] ), .op(n21648) );
  nor2_1 U25729 ( .ip1(\x[101][2] ), .ip2(n23659), .op(n21647) );
  inv_1 U25730 ( .ip(\x[101][1] ), .op(n21643) );
  nor2_1 U25731 ( .ip1(sig_in[1]), .ip2(n21643), .op(n21645) );
  inv_1 U25732 ( .ip(\x[101][0] ), .op(n21642) );
  not_ab_or_c_or_d U25733 ( .ip1(n22513), .ip2(n21643), .ip3(n23195), .ip4(
        n21642), .op(n21644) );
  not_ab_or_c_or_d U25734 ( .ip1(\x[101][2] ), .ip2(n24470), .ip3(n21645), 
        .ip4(n21644), .op(n21646) );
  not_ab_or_c_or_d U25735 ( .ip1(sig_in[3]), .ip2(n21648), .ip3(n21647), .ip4(
        n21646), .op(n21652) );
  nand2_1 U25736 ( .ip1(\x[101][5] ), .ip2(n24119), .op(n21650) );
  nand2_1 U25737 ( .ip1(\x[101][4] ), .ip2(n23721), .op(n21649) );
  nand2_1 U25738 ( .ip1(n21650), .ip2(n21649), .op(n21651) );
  not_ab_or_c_or_d U25739 ( .ip1(\x[101][3] ), .ip2(n24476), .ip3(n21652), 
        .ip4(n21651), .op(n21656) );
  nor2_1 U25740 ( .ip1(\x[101][5] ), .ip2(n24350), .op(n21655) );
  nor2_1 U25741 ( .ip1(\x[101][6] ), .ip2(n23509), .op(n21654) );
  not_ab_or_c_or_d U25742 ( .ip1(\x[101][5] ), .ip2(n23600), .ip3(\x[101][4] ), 
        .ip4(n24347), .op(n21653) );
  nor4_1 U25743 ( .ip1(n21656), .ip2(n21655), .ip3(n21654), .ip4(n21653), .op(
        n21657) );
  not_ab_or_c_or_d U25744 ( .ip1(\x[101][6] ), .ip2(n24045), .ip3(n21658), 
        .ip4(n21657), .op(n21662) );
  nor2_1 U25745 ( .ip1(\x[101][8] ), .ip2(n24358), .op(n21660) );
  nor2_1 U25746 ( .ip1(\x[101][7] ), .ip2(n24044), .op(n21659) );
  nor4_1 U25747 ( .ip1(n21662), .ip2(n21661), .ip3(n21660), .ip4(n21659), .op(
        n21663) );
  not_ab_or_c_or_d U25748 ( .ip1(\x[101][10] ), .ip2(n24370), .ip3(n21664), 
        .ip4(n21663), .op(n21665) );
  nand2_1 U25749 ( .ip1(n21666), .ip2(n21665), .op(n21672) );
  nor2_1 U25750 ( .ip1(\x[101][10] ), .ip2(n24457), .op(n21667) );
  or2_1 U25751 ( .ip1(sig_in[11]), .ip2(n21667), .op(n21670) );
  inv_1 U25752 ( .ip(\x[101][11] ), .op(n21668) );
  or2_1 U25753 ( .ip1(n21668), .ip2(n21667), .op(n21669) );
  nand2_1 U25754 ( .ip1(n21670), .ip2(n21669), .op(n21671) );
  nand2_1 U25755 ( .ip1(n21672), .ip2(n21671), .op(n21674) );
  nand2_1 U25756 ( .ip1(\x[101][11] ), .ip2(n24239), .op(n21673) );
  nand2_1 U25757 ( .ip1(n21674), .ip2(n21673), .op(n22379) );
  nand2_1 U25758 ( .ip1(\x[101][12] ), .ip2(n24233), .op(n21675) );
  nand2_1 U25759 ( .ip1(n21717), .ip2(n21675), .op(n22368) );
  nor2_1 U25760 ( .ip1(n22379), .ip2(n22368), .op(n21713) );
  nor2_1 U25761 ( .ip1(\x[100][11] ), .ip2(n24456), .op(n21677) );
  nor2_1 U25762 ( .ip1(\x[100][10] ), .ip2(n24457), .op(n21676) );
  nor2_1 U25763 ( .ip1(n21677), .ip2(n21676), .op(n21706) );
  inv_1 U25764 ( .ip(n21706), .op(n21678) );
  nand2_1 U25765 ( .ip1(\x[100][11] ), .ip2(n24239), .op(n21683) );
  nand2_1 U25766 ( .ip1(n21678), .ip2(n21683), .op(n22390) );
  nor2_1 U25767 ( .ip1(n23981), .ip2(\x[100][9] ), .op(n21705) );
  inv_1 U25768 ( .ip(n21705), .op(n21679) );
  nand3_1 U25769 ( .ip1(\x[100][8] ), .ip2(n24491), .ip3(n21679), .op(n21682)
         );
  nand2_1 U25770 ( .ip1(\x[100][9] ), .ip2(n23981), .op(n21681) );
  nand2_1 U25771 ( .ip1(\x[100][10] ), .ip2(n23146), .op(n21680) );
  nand4_1 U25772 ( .ip1(n21683), .ip2(n21682), .ip3(n21681), .ip4(n21680), 
        .op(n21684) );
  nand2_1 U25773 ( .ip1(n22390), .ip2(n21684), .op(n22386) );
  and2_1 U25774 ( .ip1(n24461), .ip2(\x[100][7] ), .op(n21701) );
  inv_1 U25775 ( .ip(\x[100][5] ), .op(n21699) );
  nor2_1 U25776 ( .ip1(sig_in[5]), .ip2(n21699), .op(n21696) );
  inv_1 U25777 ( .ip(\x[100][3] ), .op(n21694) );
  and2_1 U25778 ( .ip1(n24335), .ip2(\x[100][2] ), .op(n21691) );
  nand2_1 U25779 ( .ip1(\x[100][1] ), .ip2(n21685), .op(n21689) );
  nand2_1 U25780 ( .ip1(\x[100][0] ), .ip2(n24143), .op(n21688) );
  nor2_1 U25781 ( .ip1(\x[100][2] ), .ip2(n23659), .op(n21687) );
  nor2_1 U25782 ( .ip1(\x[100][1] ), .ip2(n20652), .op(n21686) );
  not_ab_or_c_or_d U25783 ( .ip1(n21689), .ip2(n21688), .ip3(n21687), .ip4(
        n21686), .op(n21690) );
  not_ab_or_c_or_d U25784 ( .ip1(\x[100][3] ), .ip2(n22525), .ip3(n21691), 
        .ip4(n21690), .op(n21693) );
  nor2_1 U25785 ( .ip1(\x[100][4] ), .ip2(n24256), .op(n21692) );
  not_ab_or_c_or_d U25786 ( .ip1(n24251), .ip2(n21694), .ip3(n21693), .ip4(
        n21692), .op(n21695) );
  not_ab_or_c_or_d U25787 ( .ip1(\x[100][4] ), .ip2(n24347), .ip3(n21696), 
        .ip4(n21695), .op(n21698) );
  nor2_1 U25788 ( .ip1(\x[100][6] ), .ip2(n23770), .op(n21697) );
  not_ab_or_c_or_d U25789 ( .ip1(n22833), .ip2(n21699), .ip3(n21698), .ip4(
        n21697), .op(n21700) );
  not_ab_or_c_or_d U25790 ( .ip1(\x[100][6] ), .ip2(n23770), .ip3(n21701), 
        .ip4(n21700), .op(n21704) );
  nor2_1 U25791 ( .ip1(\x[100][8] ), .ip2(n24358), .op(n21703) );
  nor2_1 U25792 ( .ip1(\x[100][7] ), .ip2(n24492), .op(n21702) );
  nor4_1 U25793 ( .ip1(n21705), .ip2(n21704), .ip3(n21703), .ip4(n21702), .op(
        n22391) );
  nand2_1 U25794 ( .ip1(n21706), .ip2(n22391), .op(n21711) );
  or2_1 U25795 ( .ip1(n24185), .ip2(\x[100][14] ), .op(n21707) );
  nand2_1 U25796 ( .ip1(n21708), .ip2(n21707), .op(n22400) );
  nor2_1 U25797 ( .ip1(\x[100][13] ), .ip2(n24376), .op(n21710) );
  nor2_1 U25798 ( .ip1(\x[100][12] ), .ip2(n24079), .op(n21709) );
  or2_1 U25799 ( .ip1(n21710), .ip2(n21709), .op(n22393) );
  not_ab_or_c_or_d U25800 ( .ip1(n22386), .ip2(n21711), .ip3(n22400), .ip4(
        n22393), .op(n21712) );
  nor2_1 U25801 ( .ip1(\x[100][15] ), .ip2(n24180), .op(n22384) );
  or4_1 U25802 ( .ip1(n22367), .ip2(n21713), .ip3(n21712), .ip4(n22384), .op(
        n21714) );
  not_ab_or_c_or_d U25803 ( .ip1(n21717), .ip2(n21716), .ip3(n21715), .ip4(
        n21714), .op(n24604) );
  nand2_1 U25804 ( .ip1(\x[102][15] ), .ip2(n24180), .op(n22371) );
  and2_1 U25805 ( .ip1(n23895), .ip2(\x[102][13] ), .op(n21719) );
  nor2_1 U25806 ( .ip1(\x[102][15] ), .ip2(n24180), .op(n21718) );
  not_ab_or_c_or_d U25807 ( .ip1(\x[102][14] ), .ip2(n24382), .ip3(n21719), 
        .ip4(n21718), .op(n22377) );
  nand2_1 U25808 ( .ip1(\x[102][12] ), .ip2(n24449), .op(n21720) );
  nand2_1 U25809 ( .ip1(n22377), .ip2(n21720), .op(n22372) );
  and2_1 U25810 ( .ip1(n24451), .ip2(\x[103][10] ), .op(n21747) );
  inv_1 U25811 ( .ip(\x[103][9] ), .op(n21745) );
  and2_1 U25812 ( .ip1(n23804), .ip2(\x[103][8] ), .op(n21742) );
  inv_1 U25813 ( .ip(\x[103][7] ), .op(n21740) );
  nor2_1 U25814 ( .ip1(n17732), .ip2(n21740), .op(n21737) );
  inv_1 U25815 ( .ip(\x[103][3] ), .op(n21727) );
  nor2_1 U25816 ( .ip1(\x[103][2] ), .ip2(n23717), .op(n21726) );
  inv_1 U25817 ( .ip(\x[103][1] ), .op(n21722) );
  nor2_1 U25818 ( .ip1(sig_in[1]), .ip2(n21722), .op(n21724) );
  inv_1 U25819 ( .ip(\x[103][0] ), .op(n21721) );
  not_ab_or_c_or_d U25820 ( .ip1(n22513), .ip2(n21722), .ip3(n23195), .ip4(
        n21721), .op(n21723) );
  not_ab_or_c_or_d U25821 ( .ip1(\x[103][2] ), .ip2(n24107), .ip3(n21724), 
        .ip4(n21723), .op(n21725) );
  not_ab_or_c_or_d U25822 ( .ip1(n24251), .ip2(n21727), .ip3(n21726), .ip4(
        n21725), .op(n21731) );
  nand2_1 U25823 ( .ip1(\x[103][5] ), .ip2(n24119), .op(n21729) );
  nand2_1 U25824 ( .ip1(\x[103][4] ), .ip2(n24256), .op(n21728) );
  nand2_1 U25825 ( .ip1(n21729), .ip2(n21728), .op(n21730) );
  not_ab_or_c_or_d U25826 ( .ip1(\x[103][3] ), .ip2(n24476), .ip3(n21731), 
        .ip4(n21730), .op(n21735) );
  nor2_1 U25827 ( .ip1(\x[103][5] ), .ip2(n24350), .op(n21734) );
  nor2_1 U25828 ( .ip1(\x[103][6] ), .ip2(n24355), .op(n21733) );
  not_ab_or_c_or_d U25829 ( .ip1(\x[103][5] ), .ip2(n24482), .ip3(\x[103][4] ), 
        .ip4(n24256), .op(n21732) );
  nor4_1 U25830 ( .ip1(n21735), .ip2(n21734), .ip3(n21733), .ip4(n21732), .op(
        n21736) );
  not_ab_or_c_or_d U25831 ( .ip1(\x[103][6] ), .ip2(n23509), .ip3(n21737), 
        .ip4(n21736), .op(n21739) );
  nor2_1 U25832 ( .ip1(\x[103][8] ), .ip2(n24358), .op(n21738) );
  not_ab_or_c_or_d U25833 ( .ip1(sig_in[7]), .ip2(n21740), .ip3(n21739), .ip4(
        n21738), .op(n21741) );
  not_ab_or_c_or_d U25834 ( .ip1(\x[103][9] ), .ip2(n23981), .ip3(n21742), 
        .ip4(n21741), .op(n21744) );
  nor2_1 U25835 ( .ip1(\x[103][10] ), .ip2(n24370), .op(n21743) );
  not_ab_or_c_or_d U25836 ( .ip1(sig_in[9]), .ip2(n21745), .ip3(n21744), .ip4(
        n21743), .op(n21746) );
  not_ab_or_c_or_d U25837 ( .ip1(\x[103][11] ), .ip2(n24239), .ip3(n21747), 
        .ip4(n21746), .op(n21749) );
  nor2_1 U25838 ( .ip1(\x[103][11] ), .ip2(n24456), .op(n21748) );
  nor2_1 U25839 ( .ip1(n21749), .ip2(n21748), .op(n22358) );
  and2_1 U25840 ( .ip1(n24332), .ip2(\x[103][13] ), .op(n21750) );
  nor2_1 U25841 ( .ip1(\x[103][15] ), .ip2(n24329), .op(n21756) );
  not_ab_or_c_or_d U25842 ( .ip1(\x[103][14] ), .ip2(n24382), .ip3(n21750), 
        .ip4(n21756), .op(n21755) );
  nand2_1 U25843 ( .ip1(\x[103][12] ), .ip2(n24450), .op(n21751) );
  nand2_1 U25844 ( .ip1(n21755), .ip2(n21751), .op(n22357) );
  nor2_1 U25845 ( .ip1(n22358), .ip2(n22357), .op(n21802) );
  nor2_1 U25846 ( .ip1(\x[103][13] ), .ip2(n24376), .op(n21753) );
  nor2_1 U25847 ( .ip1(\x[103][12] ), .ip2(n24233), .op(n21752) );
  nor2_1 U25848 ( .ip1(n21753), .ip2(n21752), .op(n22359) );
  inv_1 U25849 ( .ip(n22359), .op(n21754) );
  nand2_1 U25850 ( .ip1(n21755), .ip2(n21754), .op(n21800) );
  nor3_1 U25851 ( .ip1(n21756), .ip2(\x[103][14] ), .ip3(n24382), .op(n21757)
         );
  or2_1 U25852 ( .ip1(\x[103][15] ), .ip2(n21757), .op(n21759) );
  or2_1 U25853 ( .ip1(n24384), .ip2(n21757), .op(n21758) );
  nand2_1 U25854 ( .ip1(n21759), .ip2(n21758), .op(n22363) );
  nand2_1 U25855 ( .ip1(\x[102][10] ), .ip2(n23146), .op(n21786) );
  nor2_1 U25856 ( .ip1(\x[102][9] ), .ip2(n24269), .op(n21782) );
  inv_1 U25857 ( .ip(\x[102][8] ), .op(n21760) );
  nor3_1 U25858 ( .ip1(sig_in[8]), .ip2(n21782), .ip3(n21760), .op(n21784) );
  nor2_1 U25859 ( .ip1(\x[102][7] ), .ip2(n24044), .op(n21781) );
  nor2_1 U25860 ( .ip1(\x[102][8] ), .ip2(n24358), .op(n21780) );
  and2_1 U25861 ( .ip1(n24045), .ip2(\x[102][6] ), .op(n21774) );
  inv_1 U25862 ( .ip(\x[102][4] ), .op(n21772) );
  nor2_1 U25863 ( .ip1(n24462), .ip2(n21772), .op(n21769) );
  inv_1 U25864 ( .ip(\x[102][3] ), .op(n21767) );
  inv_1 U25865 ( .ip(\x[102][1] ), .op(n21762) );
  nor2_1 U25866 ( .ip1(sig_in[1]), .ip2(n21762), .op(n21764) );
  inv_1 U25867 ( .ip(\x[102][0] ), .op(n21761) );
  not_ab_or_c_or_d U25868 ( .ip1(n22513), .ip2(n21762), .ip3(n23195), .ip4(
        n21761), .op(n21763) );
  not_ab_or_c_or_d U25869 ( .ip1(\x[102][2] ), .ip2(n24470), .ip3(n21764), 
        .ip4(n21763), .op(n21766) );
  nor2_1 U25870 ( .ip1(\x[102][2] ), .ip2(n23659), .op(n21765) );
  not_ab_or_c_or_d U25871 ( .ip1(sig_in[3]), .ip2(n21767), .ip3(n21766), .ip4(
        n21765), .op(n21768) );
  not_ab_or_c_or_d U25872 ( .ip1(\x[102][3] ), .ip2(n24476), .ip3(n21769), 
        .ip4(n21768), .op(n21771) );
  nor2_1 U25873 ( .ip1(\x[102][5] ), .ip2(n24350), .op(n21770) );
  not_ab_or_c_or_d U25874 ( .ip1(sig_in[4]), .ip2(n21772), .ip3(n21771), .ip4(
        n21770), .op(n21773) );
  not_ab_or_c_or_d U25875 ( .ip1(\x[102][5] ), .ip2(n23600), .ip3(n21774), 
        .ip4(n21773), .op(n21776) );
  nor2_1 U25876 ( .ip1(n24045), .ip2(\x[102][6] ), .op(n21775) );
  nor2_1 U25877 ( .ip1(n21776), .ip2(n21775), .op(n21778) );
  and2_1 U25878 ( .ip1(n24461), .ip2(\x[102][7] ), .op(n21777) );
  nor2_1 U25879 ( .ip1(n21778), .ip2(n21777), .op(n21779) );
  nor4_1 U25880 ( .ip1(n21782), .ip2(n21781), .ip3(n21780), .ip4(n21779), .op(
        n21783) );
  not_ab_or_c_or_d U25881 ( .ip1(\x[102][9] ), .ip2(n24164), .ip3(n21784), 
        .ip4(n21783), .op(n21785) );
  nand2_1 U25882 ( .ip1(n21786), .ip2(n21785), .op(n21792) );
  nor2_1 U25883 ( .ip1(\x[102][10] ), .ip2(n24457), .op(n21787) );
  or2_1 U25884 ( .ip1(sig_in[11]), .ip2(n21787), .op(n21790) );
  inv_1 U25885 ( .ip(\x[102][11] ), .op(n21788) );
  or2_1 U25886 ( .ip1(n21788), .ip2(n21787), .op(n21789) );
  nand2_1 U25887 ( .ip1(n21790), .ip2(n21789), .op(n21791) );
  nand2_1 U25888 ( .ip1(n21792), .ip2(n21791), .op(n21795) );
  nand2_1 U25889 ( .ip1(\x[102][11] ), .ip2(n21793), .op(n21794) );
  nand2_1 U25890 ( .ip1(n21795), .ip2(n21794), .op(n22373) );
  inv_1 U25891 ( .ip(\x[102][14] ), .op(n21798) );
  nor2_1 U25892 ( .ip1(\x[102][12] ), .ip2(n24233), .op(n21797) );
  nor2_1 U25893 ( .ip1(\x[102][13] ), .ip2(n24376), .op(n21796) );
  not_ab_or_c_or_d U25894 ( .ip1(sig_in[14]), .ip2(n21798), .ip3(n21797), 
        .ip4(n21796), .op(n22370) );
  nand3_1 U25895 ( .ip1(n22373), .ip2(n22370), .ip3(n22371), .op(n21799) );
  nand3_1 U25896 ( .ip1(n21800), .ip2(n22363), .ip3(n21799), .op(n21801) );
  not_ab_or_c_or_d U25897 ( .ip1(n22371), .ip2(n22372), .ip3(n21802), .ip4(
        n21801), .op(n24580) );
  nand2_1 U25898 ( .ip1(\x[104][15] ), .ip2(n24329), .op(n21887) );
  and2_1 U25899 ( .ip1(n23895), .ip2(\x[104][13] ), .op(n21803) );
  nor2_1 U25900 ( .ip1(\x[104][15] ), .ip2(n24180), .op(n22348) );
  not_ab_or_c_or_d U25901 ( .ip1(\x[104][14] ), .ip2(n24382), .ip3(n21803), 
        .ip4(n22348), .op(n22355) );
  nand2_1 U25902 ( .ip1(\x[104][12] ), .ip2(n24450), .op(n22352) );
  nand2_1 U25903 ( .ip1(n22355), .ip2(n22352), .op(n21886) );
  nand2_1 U25904 ( .ip1(\x[105][8] ), .ip2(n23804), .op(n21824) );
  nor2_1 U25905 ( .ip1(\x[105][5] ), .ip2(n23283), .op(n21813) );
  inv_1 U25906 ( .ip(\x[105][4] ), .op(n21804) );
  nor3_1 U25907 ( .ip1(n24462), .ip2(n21813), .ip3(n21804), .op(n21816) );
  and2_1 U25908 ( .ip1(n24107), .ip2(\x[105][2] ), .op(n21810) );
  nand2_1 U25909 ( .ip1(\x[105][1] ), .ip2(n20652), .op(n21808) );
  nand2_1 U25910 ( .ip1(\x[105][0] ), .ip2(n24143), .op(n21807) );
  nor2_1 U25911 ( .ip1(\x[105][2] ), .ip2(n23659), .op(n21806) );
  nor2_1 U25912 ( .ip1(\x[105][1] ), .ip2(n20652), .op(n21805) );
  not_ab_or_c_or_d U25913 ( .ip1(n21808), .ip2(n21807), .ip3(n21806), .ip4(
        n21805), .op(n21809) );
  not_ab_or_c_or_d U25914 ( .ip1(\x[105][3] ), .ip2(n22525), .ip3(n21810), 
        .ip4(n21809), .op(n21814) );
  nor2_1 U25915 ( .ip1(\x[105][3] ), .ip2(n24342), .op(n21812) );
  nor2_1 U25916 ( .ip1(\x[105][4] ), .ip2(n23860), .op(n21811) );
  nor4_1 U25917 ( .ip1(n21814), .ip2(n21813), .ip3(n21812), .ip4(n21811), .op(
        n21815) );
  not_ab_or_c_or_d U25918 ( .ip1(\x[105][5] ), .ip2(n24482), .ip3(n21816), 
        .ip4(n21815), .op(n21820) );
  nand2_1 U25919 ( .ip1(\x[105][6] ), .ip2(n24485), .op(n21819) );
  nor2_1 U25920 ( .ip1(\x[105][6] ), .ip2(n24485), .op(n21818) );
  nor2_1 U25921 ( .ip1(\x[105][7] ), .ip2(n24492), .op(n21817) );
  not_ab_or_c_or_d U25922 ( .ip1(n21820), .ip2(n21819), .ip3(n21818), .ip4(
        n21817), .op(n21821) );
  or2_1 U25923 ( .ip1(\x[105][7] ), .ip2(n21821), .op(n21823) );
  or2_1 U25924 ( .ip1(n24044), .ip2(n21821), .op(n21822) );
  nand2_1 U25925 ( .ip1(n21823), .ip2(n21822), .op(n22328) );
  nand2_1 U25926 ( .ip1(n21824), .ip2(n22328), .op(n21827) );
  nor2_1 U25927 ( .ip1(\x[105][9] ), .ip2(n24043), .op(n22322) );
  or2_1 U25928 ( .ip1(n23779), .ip2(n22322), .op(n21826) );
  inv_1 U25929 ( .ip(\x[105][8] ), .op(n22323) );
  or2_1 U25930 ( .ip1(n22323), .ip2(n22322), .op(n21825) );
  nand2_1 U25931 ( .ip1(n21826), .ip2(n21825), .op(n22330) );
  nand2_1 U25932 ( .ip1(n21827), .ip2(n22330), .op(n21829) );
  and2_1 U25933 ( .ip1(n24451), .ip2(\x[105][10] ), .op(n21828) );
  and2_1 U25934 ( .ip1(n24371), .ip2(\x[105][11] ), .op(n21832) );
  not_ab_or_c_or_d U25935 ( .ip1(\x[105][9] ), .ip2(n23981), .ip3(n21828), 
        .ip4(n21832), .op(n22325) );
  nand2_1 U25936 ( .ip1(n21829), .ip2(n22325), .op(n21836) );
  nor2_1 U25937 ( .ip1(\x[105][11] ), .ip2(n24456), .op(n21831) );
  nor2_1 U25938 ( .ip1(\x[105][10] ), .ip2(n24457), .op(n21830) );
  nor2_1 U25939 ( .ip1(n21831), .ip2(n21830), .op(n22331) );
  or2_1 U25940 ( .ip1(n21832), .ip2(n22331), .op(n22327) );
  nand2_1 U25941 ( .ip1(\x[105][13] ), .ip2(n24235), .op(n21834) );
  nand2_1 U25942 ( .ip1(\x[105][12] ), .ip2(n24450), .op(n21833) );
  nand2_1 U25943 ( .ip1(n21834), .ip2(n21833), .op(n22337) );
  nand2_1 U25944 ( .ip1(\x[105][14] ), .ip2(n24230), .op(n21835) );
  nor2_1 U25945 ( .ip1(n24384), .ip2(\x[105][15] ), .op(n21875) );
  inv_1 U25946 ( .ip(n21875), .op(n22345) );
  nand2_1 U25947 ( .ip1(n21835), .ip2(n22345), .op(n21880) );
  not_ab_or_c_or_d U25948 ( .ip1(n21836), .ip2(n22327), .ip3(n22337), .ip4(
        n21880), .op(n21885) );
  inv_1 U25949 ( .ip(\x[104][11] ), .op(n21867) );
  and2_1 U25950 ( .ip1(n24451), .ip2(\x[104][10] ), .op(n21864) );
  inv_1 U25951 ( .ip(\x[104][9] ), .op(n21862) );
  and2_1 U25952 ( .ip1(n23804), .ip2(\x[104][8] ), .op(n21859) );
  nor2_1 U25953 ( .ip1(n23600), .ip2(\x[104][5] ), .op(n21852) );
  and2_1 U25954 ( .ip1(n23860), .ip2(\x[104][4] ), .op(n21850) );
  inv_1 U25955 ( .ip(\x[104][3] ), .op(n21848) );
  inv_1 U25956 ( .ip(\x[104][1] ), .op(n21838) );
  nor2_1 U25957 ( .ip1(sig_in[1]), .ip2(n21838), .op(n21840) );
  inv_1 U25958 ( .ip(\x[104][0] ), .op(n21837) );
  not_ab_or_c_or_d U25959 ( .ip1(n22513), .ip2(n21838), .ip3(n23195), .ip4(
        n21837), .op(n21839) );
  not_ab_or_c_or_d U25960 ( .ip1(\x[104][2] ), .ip2(n24107), .ip3(n21840), 
        .ip4(n21839), .op(n21842) );
  nor2_1 U25961 ( .ip1(\x[104][2] ), .ip2(n23659), .op(n21841) );
  nor2_1 U25962 ( .ip1(n21842), .ip2(n21841), .op(n21843) );
  or2_1 U25963 ( .ip1(\x[104][3] ), .ip2(n21843), .op(n21845) );
  or2_1 U25964 ( .ip1(n22525), .ip2(n21843), .op(n21844) );
  nand2_1 U25965 ( .ip1(n21845), .ip2(n21844), .op(n21847) );
  nor2_1 U25966 ( .ip1(\x[104][4] ), .ip2(n24347), .op(n21846) );
  not_ab_or_c_or_d U25967 ( .ip1(n23251), .ip2(n21848), .ip3(n21847), .ip4(
        n21846), .op(n21849) );
  not_ab_or_c_or_d U25968 ( .ip1(\x[104][5] ), .ip2(n24482), .ip3(n21850), 
        .ip4(n21849), .op(n21851) );
  or2_1 U25969 ( .ip1(n21852), .ip2(n21851), .op(n21855) );
  nor2_1 U25970 ( .ip1(\x[104][7] ), .ip2(n24044), .op(n21854) );
  nor3_1 U25971 ( .ip1(sig_in[6]), .ip2(n21855), .ip3(n21854), .op(n21857) );
  inv_1 U25972 ( .ip(\x[104][6] ), .op(n21853) );
  not_ab_or_c_or_d U25973 ( .ip1(n21855), .ip2(sig_in[6]), .ip3(n21854), .ip4(
        n21853), .op(n21856) );
  or2_1 U25974 ( .ip1(n21857), .ip2(n21856), .op(n21858) );
  not_ab_or_c_or_d U25975 ( .ip1(\x[104][7] ), .ip2(n24142), .ip3(n21859), 
        .ip4(n21858), .op(n21861) );
  nor2_1 U25976 ( .ip1(\x[104][8] ), .ip2(n24100), .op(n21860) );
  not_ab_or_c_or_d U25977 ( .ip1(sig_in[9]), .ip2(n21862), .ip3(n21861), .ip4(
        n21860), .op(n21863) );
  not_ab_or_c_or_d U25978 ( .ip1(\x[104][9] ), .ip2(n24164), .ip3(n21864), 
        .ip4(n21863), .op(n21866) );
  nor2_1 U25979 ( .ip1(\x[104][10] ), .ip2(n24457), .op(n21865) );
  not_ab_or_c_or_d U25980 ( .ip1(sig_in[11]), .ip2(n21867), .ip3(n21866), 
        .ip4(n21865), .op(n21868) );
  or2_1 U25981 ( .ip1(\x[104][11] ), .ip2(n21868), .op(n21870) );
  or2_1 U25982 ( .ip1(n24371), .ip2(n21868), .op(n21869) );
  nand2_1 U25983 ( .ip1(n21870), .ip2(n21869), .op(n22351) );
  or2_1 U25984 ( .ip1(n24382), .ip2(\x[104][14] ), .op(n21871) );
  nand2_1 U25985 ( .ip1(n21887), .ip2(n21871), .op(n22350) );
  nor2_1 U25986 ( .ip1(\x[104][13] ), .ip2(n24376), .op(n21873) );
  nor2_1 U25987 ( .ip1(\x[104][12] ), .ip2(n24233), .op(n21872) );
  nor2_1 U25988 ( .ip1(n21873), .ip2(n21872), .op(n22353) );
  inv_1 U25989 ( .ip(n22353), .op(n21874) );
  nor3_1 U25990 ( .ip1(n22351), .ip2(n22350), .ip3(n21874), .op(n21883) );
  and2_1 U25991 ( .ip1(n24186), .ip2(\x[105][15] ), .op(n22340) );
  nor3_1 U25992 ( .ip1(\x[105][14] ), .ip2(n21875), .ip3(n24185), .op(n21882)
         );
  nor2_1 U25993 ( .ip1(\x[105][13] ), .ip2(n24376), .op(n21876) );
  or2_1 U25994 ( .ip1(n17845), .ip2(n21876), .op(n21879) );
  inv_1 U25995 ( .ip(\x[105][12] ), .op(n21877) );
  or2_1 U25996 ( .ip1(n21877), .ip2(n21876), .op(n21878) );
  nand2_1 U25997 ( .ip1(n21879), .ip2(n21878), .op(n22332) );
  nor2_1 U25998 ( .ip1(n22332), .ip2(n21880), .op(n21881) );
  or4_1 U25999 ( .ip1(n21883), .ip2(n22340), .ip3(n21882), .ip4(n21881), .op(
        n21884) );
  not_ab_or_c_or_d U26000 ( .ip1(n21887), .ip2(n21886), .ip3(n21885), .ip4(
        n21884), .op(n24589) );
  nand2_1 U26001 ( .ip1(\x[106][15] ), .ip2(n24180), .op(n21982) );
  or2_1 U26002 ( .ip1(n24329), .ip2(\x[106][15] ), .op(n22343) );
  nand2_1 U26003 ( .ip1(\x[106][14] ), .ip2(n23938), .op(n21888) );
  nand2_1 U26004 ( .ip1(n22343), .ip2(n21888), .op(n22319) );
  and2_1 U26005 ( .ip1(\x[106][11] ), .ip2(n24239), .op(n21891) );
  nor2_1 U26006 ( .ip1(\x[106][11] ), .ip2(n24456), .op(n21890) );
  nor2_1 U26007 ( .ip1(\x[106][10] ), .ip2(n24457), .op(n21889) );
  nor2_1 U26008 ( .ip1(n21890), .ip2(n21889), .op(n21924) );
  or2_1 U26009 ( .ip1(n21891), .ip2(n21924), .op(n22321) );
  and2_1 U26010 ( .ip1(n24451), .ip2(\x[106][10] ), .op(n21892) );
  not_ab_or_c_or_d U26011 ( .ip1(\x[106][9] ), .ip2(n24269), .ip3(n21892), 
        .ip4(n21891), .op(n22316) );
  inv_1 U26012 ( .ip(\x[106][8] ), .op(n21921) );
  nor2_1 U26013 ( .ip1(n24164), .ip2(\x[106][9] ), .op(n21920) );
  or3_1 U26014 ( .ip1(n23779), .ip2(n21921), .ip3(n21920), .op(n21893) );
  nand2_1 U26015 ( .ip1(n22316), .ip2(n21893), .op(n21894) );
  nand2_1 U26016 ( .ip1(n22321), .ip2(n21894), .op(n21929) );
  inv_1 U26017 ( .ip(\x[106][7] ), .op(n21917) );
  nor2_1 U26018 ( .ip1(n17732), .ip2(n21917), .op(n21915) );
  inv_1 U26019 ( .ip(\x[106][5] ), .op(n21913) );
  inv_1 U26020 ( .ip(\x[106][4] ), .op(n21905) );
  nor2_1 U26021 ( .ip1(n24462), .ip2(n21905), .op(n21903) );
  inv_1 U26022 ( .ip(\x[106][3] ), .op(n21901) );
  inv_1 U26023 ( .ip(\x[106][1] ), .op(n21896) );
  nor2_1 U26024 ( .ip1(sig_in[1]), .ip2(n21896), .op(n21898) );
  inv_1 U26025 ( .ip(\x[106][0] ), .op(n21895) );
  not_ab_or_c_or_d U26026 ( .ip1(n22513), .ip2(n21896), .ip3(n23195), .ip4(
        n21895), .op(n21897) );
  not_ab_or_c_or_d U26027 ( .ip1(\x[106][2] ), .ip2(n24470), .ip3(n21898), 
        .ip4(n21897), .op(n21900) );
  nor2_1 U26028 ( .ip1(\x[106][2] ), .ip2(n23659), .op(n21899) );
  not_ab_or_c_or_d U26029 ( .ip1(n24251), .ip2(n21901), .ip3(n21900), .ip4(
        n21899), .op(n21902) );
  not_ab_or_c_or_d U26030 ( .ip1(\x[106][3] ), .ip2(n22525), .ip3(n21903), 
        .ip4(n21902), .op(n21904) );
  or2_1 U26031 ( .ip1(sig_in[4]), .ip2(n21904), .op(n21907) );
  or2_1 U26032 ( .ip1(n21905), .ip2(n21904), .op(n21906) );
  nand2_1 U26033 ( .ip1(n21907), .ip2(n21906), .op(n21908) );
  or2_1 U26034 ( .ip1(\x[106][5] ), .ip2(n21908), .op(n21910) );
  or2_1 U26035 ( .ip1(n24482), .ip2(n21908), .op(n21909) );
  nand2_1 U26036 ( .ip1(n21910), .ip2(n21909), .op(n21912) );
  nor2_1 U26037 ( .ip1(\x[106][6] ), .ip2(n24485), .op(n21911) );
  not_ab_or_c_or_d U26038 ( .ip1(n22833), .ip2(n21913), .ip3(n21912), .ip4(
        n21911), .op(n21914) );
  not_ab_or_c_or_d U26039 ( .ip1(\x[106][6] ), .ip2(n24045), .ip3(n21915), 
        .ip4(n21914), .op(n21916) );
  or2_1 U26040 ( .ip1(sig_in[7]), .ip2(n21916), .op(n21919) );
  or2_1 U26041 ( .ip1(n21917), .ip2(n21916), .op(n21918) );
  nand2_1 U26042 ( .ip1(n21919), .ip2(n21918), .op(n22311) );
  or2_1 U26043 ( .ip1(n23779), .ip2(n21920), .op(n21923) );
  or2_1 U26044 ( .ip1(n21921), .ip2(n21920), .op(n21922) );
  nand2_1 U26045 ( .ip1(n21923), .ip2(n21922), .op(n22314) );
  nand3_1 U26046 ( .ip1(n21924), .ip2(n22311), .ip3(n22314), .op(n21928) );
  or2_1 U26047 ( .ip1(n24382), .ip2(\x[106][14] ), .op(n21925) );
  nand2_1 U26048 ( .ip1(n21925), .ip2(n21982), .op(n22344) );
  nor2_1 U26049 ( .ip1(\x[106][13] ), .ip2(n24376), .op(n21927) );
  nor2_1 U26050 ( .ip1(\x[106][12] ), .ip2(n24233), .op(n21926) );
  or2_1 U26051 ( .ip1(n21927), .ip2(n21926), .op(n22309) );
  not_ab_or_c_or_d U26052 ( .ip1(n21929), .ip2(n21928), .ip3(n22344), .ip4(
        n22309), .op(n21981) );
  nand2_1 U26053 ( .ip1(\x[107][14] ), .ip2(n24327), .op(n21969) );
  and2_1 U26054 ( .ip1(n24332), .ip2(\x[107][13] ), .op(n21963) );
  inv_1 U26055 ( .ip(\x[107][11] ), .op(n21961) );
  nor2_1 U26056 ( .ip1(\x[107][10] ), .ip2(n24457), .op(n21960) );
  and2_1 U26057 ( .ip1(n23804), .ip2(\x[107][8] ), .op(n21953) );
  inv_1 U26058 ( .ip(\x[107][7] ), .op(n21951) );
  nor2_1 U26059 ( .ip1(sig_in[7]), .ip2(n21951), .op(n21948) );
  inv_1 U26060 ( .ip(\x[107][5] ), .op(n21946) );
  nor2_1 U26061 ( .ip1(sig_in[5]), .ip2(n21946), .op(n21943) );
  inv_1 U26062 ( .ip(\x[107][3] ), .op(n21941) );
  and2_1 U26063 ( .ip1(n24335), .ip2(\x[107][2] ), .op(n21938) );
  inv_1 U26064 ( .ip(\x[107][1] ), .op(n21931) );
  inv_1 U26065 ( .ip(\x[107][0] ), .op(n21930) );
  not_ab_or_c_or_d U26066 ( .ip1(n22513), .ip2(n21931), .ip3(n23195), .ip4(
        n21930), .op(n21932) );
  or2_1 U26067 ( .ip1(\x[107][1] ), .ip2(n21932), .op(n21934) );
  or2_1 U26068 ( .ip1(n20652), .ip2(n21932), .op(n21933) );
  nand2_1 U26069 ( .ip1(n21934), .ip2(n21933), .op(n21936) );
  nor2_1 U26070 ( .ip1(\x[107][2] ), .ip2(n23659), .op(n21935) );
  nor2_1 U26071 ( .ip1(n21936), .ip2(n21935), .op(n21937) );
  not_ab_or_c_or_d U26072 ( .ip1(\x[107][3] ), .ip2(n24476), .ip3(n21938), 
        .ip4(n21937), .op(n21940) );
  nor2_1 U26073 ( .ip1(\x[107][4] ), .ip2(n23721), .op(n21939) );
  not_ab_or_c_or_d U26074 ( .ip1(n23251), .ip2(n21941), .ip3(n21940), .ip4(
        n21939), .op(n21942) );
  not_ab_or_c_or_d U26075 ( .ip1(\x[107][4] ), .ip2(n24347), .ip3(n21943), 
        .ip4(n21942), .op(n21945) );
  nor2_1 U26076 ( .ip1(\x[107][6] ), .ip2(n23509), .op(n21944) );
  not_ab_or_c_or_d U26077 ( .ip1(n22833), .ip2(n21946), .ip3(n21945), .ip4(
        n21944), .op(n21947) );
  not_ab_or_c_or_d U26078 ( .ip1(\x[107][6] ), .ip2(n24485), .ip3(n21948), 
        .ip4(n21947), .op(n21950) );
  nor2_1 U26079 ( .ip1(\x[107][8] ), .ip2(n24100), .op(n21949) );
  not_ab_or_c_or_d U26080 ( .ip1(sig_in[7]), .ip2(n21951), .ip3(n21950), .ip4(
        n21949), .op(n21952) );
  not_ab_or_c_or_d U26081 ( .ip1(\x[107][9] ), .ip2(n24043), .ip3(n21953), 
        .ip4(n21952), .op(n21955) );
  nor2_1 U26082 ( .ip1(\x[107][9] ), .ip2(n24455), .op(n21954) );
  nor2_1 U26083 ( .ip1(n21955), .ip2(n21954), .op(n21956) );
  or2_1 U26084 ( .ip1(\x[107][10] ), .ip2(n21956), .op(n21958) );
  or2_1 U26085 ( .ip1(n24370), .ip2(n21956), .op(n21957) );
  nand2_1 U26086 ( .ip1(n21958), .ip2(n21957), .op(n21959) );
  not_ab_or_c_or_d U26087 ( .ip1(sig_in[11]), .ip2(n21961), .ip3(n21960), 
        .ip4(n21959), .op(n21962) );
  not_ab_or_c_or_d U26088 ( .ip1(\x[107][11] ), .ip2(n21793), .ip3(n21963), 
        .ip4(n21962), .op(n21967) );
  nor2_1 U26089 ( .ip1(n17845), .ip2(n21967), .op(n21964) );
  nor2_1 U26090 ( .ip1(\x[107][12] ), .ip2(n21964), .op(n21966) );
  nor2_1 U26091 ( .ip1(\x[107][13] ), .ip2(n24376), .op(n21965) );
  ab_or_c_or_d U26092 ( .ip1(n21967), .ip2(n17845), .ip3(n21966), .ip4(n21965), 
        .op(n21968) );
  nand2_1 U26093 ( .ip1(n21969), .ip2(n21968), .op(n22304) );
  nor2_1 U26094 ( .ip1(\x[107][14] ), .ip2(n24327), .op(n21970) );
  or2_1 U26095 ( .ip1(\x[107][15] ), .ip2(n21970), .op(n21972) );
  or2_1 U26096 ( .ip1(n24329), .ip2(n21970), .op(n21971) );
  nand2_1 U26097 ( .ip1(n21972), .ip2(n21971), .op(n22303) );
  nand2_1 U26098 ( .ip1(n22304), .ip2(n22303), .op(n21974) );
  nor2_1 U26099 ( .ip1(n24384), .ip2(\x[107][15] ), .op(n22308) );
  inv_1 U26100 ( .ip(n22308), .op(n21973) );
  nand2_1 U26101 ( .ip1(n21974), .ip2(n21973), .op(n21979) );
  inv_1 U26102 ( .ip(n22344), .op(n21977) );
  nand2_1 U26103 ( .ip1(\x[106][13] ), .ip2(n24081), .op(n21976) );
  nand2_1 U26104 ( .ip1(\x[106][12] ), .ip2(n24079), .op(n21975) );
  nand2_1 U26105 ( .ip1(n21976), .ip2(n21975), .op(n22318) );
  nand2_1 U26106 ( .ip1(n21977), .ip2(n22318), .op(n21978) );
  nand2_1 U26107 ( .ip1(n21979), .ip2(n21978), .op(n21980) );
  not_ab_or_c_or_d U26108 ( .ip1(n21982), .ip2(n22319), .ip3(n21981), .ip4(
        n21980), .op(n24524) );
  nand2_1 U26109 ( .ip1(\x[108][15] ), .ip2(n24180), .op(n22076) );
  and2_1 U26110 ( .ip1(n23895), .ip2(\x[108][13] ), .op(n21983) );
  nor2_1 U26111 ( .ip1(\x[108][15] ), .ip2(n24180), .op(n22301) );
  not_ab_or_c_or_d U26112 ( .ip1(\x[108][14] ), .ip2(n23938), .ip3(n21983), 
        .ip4(n22301), .op(n22292) );
  nand2_1 U26113 ( .ip1(\x[108][12] ), .ip2(n24233), .op(n22294) );
  nand2_1 U26114 ( .ip1(n22292), .ip2(n22294), .op(n22075) );
  nand2_1 U26115 ( .ip1(\x[108][9] ), .ip2(n24269), .op(n21986) );
  nor2_1 U26116 ( .ip1(\x[108][11] ), .ip2(n21793), .op(n21985) );
  nor2_1 U26117 ( .ip1(\x[108][10] ), .ip2(n24457), .op(n21984) );
  or2_1 U26118 ( .ip1(n21985), .ip2(n21984), .op(n21990) );
  or2_1 U26119 ( .ip1(n21986), .ip2(n21990), .op(n21989) );
  nand2_1 U26120 ( .ip1(\x[108][10] ), .ip2(n23146), .op(n21987) );
  or2_1 U26121 ( .ip1(n21987), .ip2(n21990), .op(n21988) );
  nand2_1 U26122 ( .ip1(n21989), .ip2(n21988), .op(n22016) );
  nor2_1 U26123 ( .ip1(n23981), .ip2(\x[108][9] ), .op(n21991) );
  nor2_1 U26124 ( .ip1(n21991), .ip2(n21990), .op(n22012) );
  inv_1 U26125 ( .ip(\x[108][7] ), .op(n22010) );
  nor2_1 U26126 ( .ip1(n17732), .ip2(n22010), .op(n22007) );
  inv_1 U26127 ( .ip(\x[108][5] ), .op(n22005) );
  nor2_1 U26128 ( .ip1(n22833), .ip2(n22005), .op(n22002) );
  inv_1 U26129 ( .ip(\x[108][3] ), .op(n22000) );
  and2_1 U26130 ( .ip1(n24335), .ip2(\x[108][2] ), .op(n21997) );
  nand2_1 U26131 ( .ip1(\x[108][1] ), .ip2(n21685), .op(n21995) );
  nand2_1 U26132 ( .ip1(\x[108][0] ), .ip2(n24143), .op(n21994) );
  nor2_1 U26133 ( .ip1(\x[108][2] ), .ip2(n23659), .op(n21993) );
  nor2_1 U26134 ( .ip1(\x[108][1] ), .ip2(n20652), .op(n21992) );
  not_ab_or_c_or_d U26135 ( .ip1(n21995), .ip2(n21994), .ip3(n21993), .ip4(
        n21992), .op(n21996) );
  not_ab_or_c_or_d U26136 ( .ip1(\x[108][3] ), .ip2(n22525), .ip3(n21997), 
        .ip4(n21996), .op(n21999) );
  nor2_1 U26137 ( .ip1(\x[108][4] ), .ip2(n24256), .op(n21998) );
  not_ab_or_c_or_d U26138 ( .ip1(n23251), .ip2(n22000), .ip3(n21999), .ip4(
        n21998), .op(n22001) );
  not_ab_or_c_or_d U26139 ( .ip1(\x[108][4] ), .ip2(n24347), .ip3(n22002), 
        .ip4(n22001), .op(n22004) );
  nor2_1 U26140 ( .ip1(\x[108][6] ), .ip2(n24485), .op(n22003) );
  not_ab_or_c_or_d U26141 ( .ip1(sig_in[5]), .ip2(n22005), .ip3(n22004), .ip4(
        n22003), .op(n22006) );
  not_ab_or_c_or_d U26142 ( .ip1(\x[108][6] ), .ip2(n23509), .ip3(n22007), 
        .ip4(n22006), .op(n22009) );
  nor2_1 U26143 ( .ip1(\x[108][8] ), .ip2(n24358), .op(n22008) );
  not_ab_or_c_or_d U26144 ( .ip1(sig_in[7]), .ip2(n22010), .ip3(n22009), .ip4(
        n22008), .op(n22011) );
  nand2_1 U26145 ( .ip1(n22012), .ip2(n22011), .op(n22014) );
  nand3_1 U26146 ( .ip1(n22012), .ip2(n23971), .ip3(\x[108][8] ), .op(n22013)
         );
  nand2_1 U26147 ( .ip1(n22014), .ip2(n22013), .op(n22015) );
  not_ab_or_c_or_d U26148 ( .ip1(\x[108][11] ), .ip2(n24456), .ip3(n22016), 
        .ip4(n22015), .op(n22295) );
  or2_1 U26149 ( .ip1(n24382), .ip2(\x[108][14] ), .op(n22017) );
  nand2_1 U26150 ( .ip1(n22017), .ip2(n22076), .op(n22300) );
  nor2_1 U26151 ( .ip1(\x[108][13] ), .ip2(n24137), .op(n22019) );
  nor2_1 U26152 ( .ip1(\x[108][12] ), .ip2(n24449), .op(n22018) );
  nor2_1 U26153 ( .ip1(n22019), .ip2(n22018), .op(n22293) );
  inv_1 U26154 ( .ip(n22293), .op(n22020) );
  nor3_1 U26155 ( .ip1(n22295), .ip2(n22300), .ip3(n22020), .op(n22074) );
  nand2_1 U26156 ( .ip1(n24332), .ip2(\x[109][13] ), .op(n22022) );
  nand2_1 U26157 ( .ip1(\x[109][12] ), .ip2(n24233), .op(n22021) );
  nand2_1 U26158 ( .ip1(n22022), .ip2(n22021), .op(n22283) );
  nor2_1 U26159 ( .ip1(n24239), .ip2(\x[109][11] ), .op(n22060) );
  inv_1 U26160 ( .ip(\x[109][9] ), .op(n22056) );
  and2_1 U26161 ( .ip1(n23804), .ip2(\x[109][8] ), .op(n22053) );
  inv_1 U26162 ( .ip(\x[109][6] ), .op(n22046) );
  inv_1 U26163 ( .ip(\x[109][5] ), .op(n22038) );
  nor2_1 U26164 ( .ip1(n22833), .ip2(n22038), .op(n22036) );
  inv_1 U26165 ( .ip(\x[109][3] ), .op(n22034) );
  inv_1 U26166 ( .ip(\x[109][1] ), .op(n22024) );
  nor2_1 U26167 ( .ip1(sig_in[1]), .ip2(n22024), .op(n22026) );
  inv_1 U26168 ( .ip(\x[109][0] ), .op(n22023) );
  not_ab_or_c_or_d U26169 ( .ip1(n22513), .ip2(n22024), .ip3(n23195), .ip4(
        n22023), .op(n22025) );
  not_ab_or_c_or_d U26170 ( .ip1(\x[109][2] ), .ip2(n24107), .ip3(n22026), 
        .ip4(n22025), .op(n22028) );
  nor2_1 U26171 ( .ip1(\x[109][2] ), .ip2(n23659), .op(n22027) );
  nor2_1 U26172 ( .ip1(n22028), .ip2(n22027), .op(n22029) );
  or2_1 U26173 ( .ip1(\x[109][3] ), .ip2(n22029), .op(n22031) );
  or2_1 U26174 ( .ip1(n24476), .ip2(n22029), .op(n22030) );
  nand2_1 U26175 ( .ip1(n22031), .ip2(n22030), .op(n22033) );
  nor2_1 U26176 ( .ip1(\x[109][4] ), .ip2(n23860), .op(n22032) );
  not_ab_or_c_or_d U26177 ( .ip1(n24251), .ip2(n22034), .ip3(n22033), .ip4(
        n22032), .op(n22035) );
  not_ab_or_c_or_d U26178 ( .ip1(\x[109][4] ), .ip2(n23860), .ip3(n22036), 
        .ip4(n22035), .op(n22037) );
  or2_1 U26179 ( .ip1(sig_in[5]), .ip2(n22037), .op(n22040) );
  or2_1 U26180 ( .ip1(n22038), .ip2(n22037), .op(n22039) );
  nand2_1 U26181 ( .ip1(n22040), .ip2(n22039), .op(n22041) );
  or2_1 U26182 ( .ip1(\x[109][6] ), .ip2(n22041), .op(n22043) );
  or2_1 U26183 ( .ip1(n24485), .ip2(n22041), .op(n22042) );
  nand2_1 U26184 ( .ip1(n22043), .ip2(n22042), .op(n22045) );
  nor2_1 U26185 ( .ip1(\x[109][7] ), .ip2(n24044), .op(n22044) );
  not_ab_or_c_or_d U26186 ( .ip1(sig_in[6]), .ip2(n22046), .ip3(n22045), .ip4(
        n22044), .op(n22047) );
  or2_1 U26187 ( .ip1(\x[109][7] ), .ip2(n22047), .op(n22049) );
  or2_1 U26188 ( .ip1(n24492), .ip2(n22047), .op(n22048) );
  nand2_1 U26189 ( .ip1(n22049), .ip2(n22048), .op(n22051) );
  nor2_1 U26190 ( .ip1(\x[109][8] ), .ip2(n24358), .op(n22050) );
  nor2_1 U26191 ( .ip1(n22051), .ip2(n22050), .op(n22052) );
  not_ab_or_c_or_d U26192 ( .ip1(\x[109][9] ), .ip2(n24455), .ip3(n22053), 
        .ip4(n22052), .op(n22055) );
  nor2_1 U26193 ( .ip1(\x[109][10] ), .ip2(n24457), .op(n22054) );
  not_ab_or_c_or_d U26194 ( .ip1(sig_in[9]), .ip2(n22056), .ip3(n22055), .ip4(
        n22054), .op(n22058) );
  and2_1 U26195 ( .ip1(n24451), .ip2(\x[109][10] ), .op(n22057) );
  not_ab_or_c_or_d U26196 ( .ip1(\x[109][11] ), .ip2(n24371), .ip3(n22058), 
        .ip4(n22057), .op(n22059) );
  nor2_1 U26197 ( .ip1(n22060), .ip2(n22059), .op(n22282) );
  or2_1 U26198 ( .ip1(n22283), .ip2(n22282), .op(n22065) );
  nor2_1 U26199 ( .ip1(\x[109][13] ), .ip2(n24137), .op(n22061) );
  or2_1 U26200 ( .ip1(n17845), .ip2(n22061), .op(n22064) );
  inv_1 U26201 ( .ip(\x[109][12] ), .op(n22062) );
  or2_1 U26202 ( .ip1(n22062), .ip2(n22061), .op(n22063) );
  nand2_1 U26203 ( .ip1(n22064), .ip2(n22063), .op(n22281) );
  nand2_1 U26204 ( .ip1(n22065), .ip2(n22281), .op(n22068) );
  nor2_1 U26205 ( .ip1(\x[109][15] ), .ip2(n24329), .op(n22070) );
  or2_1 U26206 ( .ip1(\x[109][14] ), .ip2(n22070), .op(n22067) );
  or2_1 U26207 ( .ip1(n24327), .ip2(n22070), .op(n22066) );
  nand2_1 U26208 ( .ip1(n22067), .ip2(n22066), .op(n22285) );
  nand2_1 U26209 ( .ip1(n22068), .ip2(n22285), .op(n22072) );
  nand2_1 U26210 ( .ip1(\x[109][15] ), .ip2(n24329), .op(n22287) );
  or2_1 U26211 ( .ip1(n24382), .ip2(\x[109][14] ), .op(n22069) );
  and2_1 U26212 ( .ip1(n22287), .ip2(n22069), .op(n22284) );
  or2_1 U26213 ( .ip1(n22284), .ip2(n22070), .op(n22071) );
  nand2_1 U26214 ( .ip1(n22072), .ip2(n22071), .op(n22073) );
  not_ab_or_c_or_d U26215 ( .ip1(n22076), .ip2(n22075), .ip3(n22074), .ip4(
        n22073), .op(n24960) );
  nand2_1 U26216 ( .ip1(\x[110][15] ), .ip2(n24329), .op(n22169) );
  and2_1 U26217 ( .ip1(n23895), .ip2(\x[110][13] ), .op(n22077) );
  nor2_1 U26218 ( .ip1(\x[110][15] ), .ip2(n24329), .op(n22275) );
  not_ab_or_c_or_d U26219 ( .ip1(\x[110][14] ), .ip2(n24327), .ip3(n22077), 
        .ip4(n22275), .op(n22272) );
  nand2_1 U26220 ( .ip1(\x[110][12] ), .ip2(n24450), .op(n22078) );
  nand2_1 U26221 ( .ip1(n22272), .ip2(n22078), .op(n22271) );
  nor2_1 U26222 ( .ip1(\x[111][13] ), .ip2(n24137), .op(n22079) );
  or2_1 U26223 ( .ip1(n17845), .ip2(n22079), .op(n22082) );
  inv_1 U26224 ( .ip(\x[111][12] ), .op(n22080) );
  or2_1 U26225 ( .ip1(n22080), .ip2(n22079), .op(n22081) );
  nand2_1 U26226 ( .ip1(n22082), .ip2(n22081), .op(n22176) );
  nor2_1 U26227 ( .ip1(\x[111][15] ), .ip2(n24180), .op(n22174) );
  or2_1 U26228 ( .ip1(n22176), .ip2(n22174), .op(n22126) );
  nor2_1 U26229 ( .ip1(\x[111][14] ), .ip2(n24327), .op(n22083) );
  or2_1 U26230 ( .ip1(\x[111][15] ), .ip2(n22083), .op(n22085) );
  or2_1 U26231 ( .ip1(n24384), .ip2(n22083), .op(n22084) );
  nand2_1 U26232 ( .ip1(n22085), .ip2(n22084), .op(n22123) );
  inv_1 U26233 ( .ip(\x[111][11] ), .op(n22115) );
  nor2_1 U26234 ( .ip1(n22115), .ip2(n17981), .op(n22117) );
  and2_1 U26235 ( .ip1(n24451), .ip2(\x[111][10] ), .op(n22112) );
  inv_1 U26236 ( .ip(\x[111][7] ), .op(n22105) );
  nor2_1 U26237 ( .ip1(n17732), .ip2(n22105), .op(n22102) );
  inv_1 U26238 ( .ip(\x[111][3] ), .op(n22092) );
  inv_1 U26239 ( .ip(\x[111][1] ), .op(n22087) );
  nor2_1 U26240 ( .ip1(sig_in[1]), .ip2(n22087), .op(n22089) );
  inv_1 U26241 ( .ip(\x[111][0] ), .op(n22086) );
  not_ab_or_c_or_d U26242 ( .ip1(n24467), .ip2(n22087), .ip3(n23195), .ip4(
        n22086), .op(n22088) );
  not_ab_or_c_or_d U26243 ( .ip1(\x[111][2] ), .ip2(n24470), .ip3(n22089), 
        .ip4(n22088), .op(n22091) );
  nor2_1 U26244 ( .ip1(\x[111][2] ), .ip2(n23659), .op(n22090) );
  not_ab_or_c_or_d U26245 ( .ip1(n24251), .ip2(n22092), .ip3(n22091), .ip4(
        n22090), .op(n22096) );
  nand2_1 U26246 ( .ip1(\x[111][5] ), .ip2(n24119), .op(n22094) );
  nand2_1 U26247 ( .ip1(\x[111][4] ), .ip2(n23721), .op(n22093) );
  nand2_1 U26248 ( .ip1(n22094), .ip2(n22093), .op(n22095) );
  not_ab_or_c_or_d U26249 ( .ip1(\x[111][3] ), .ip2(n22525), .ip3(n22096), 
        .ip4(n22095), .op(n22100) );
  nor2_1 U26250 ( .ip1(\x[111][6] ), .ip2(n24355), .op(n22099) );
  nor2_1 U26251 ( .ip1(\x[111][5] ), .ip2(n24350), .op(n22098) );
  not_ab_or_c_or_d U26252 ( .ip1(\x[111][5] ), .ip2(n23600), .ip3(\x[111][4] ), 
        .ip4(n24256), .op(n22097) );
  nor4_1 U26253 ( .ip1(n22100), .ip2(n22099), .ip3(n22098), .ip4(n22097), .op(
        n22101) );
  not_ab_or_c_or_d U26254 ( .ip1(\x[111][6] ), .ip2(n23770), .ip3(n22102), 
        .ip4(n22101), .op(n22104) );
  nor2_1 U26255 ( .ip1(\x[111][8] ), .ip2(n24358), .op(n22103) );
  not_ab_or_c_or_d U26256 ( .ip1(sig_in[7]), .ip2(n22105), .ip3(n22104), .ip4(
        n22103), .op(n22106) );
  or2_1 U26257 ( .ip1(\x[111][8] ), .ip2(n22106), .op(n22108) );
  or2_1 U26258 ( .ip1(n24100), .ip2(n22106), .op(n22107) );
  nand2_1 U26259 ( .ip1(n22108), .ip2(n22107), .op(n22110) );
  nor2_1 U26260 ( .ip1(\x[111][9] ), .ip2(n23981), .op(n22109) );
  nor2_1 U26261 ( .ip1(n22110), .ip2(n22109), .op(n22111) );
  not_ab_or_c_or_d U26262 ( .ip1(\x[111][9] ), .ip2(n24455), .ip3(n22112), 
        .ip4(n22111), .op(n22114) );
  nor2_1 U26263 ( .ip1(\x[111][10] ), .ip2(n24457), .op(n22113) );
  not_ab_or_c_or_d U26264 ( .ip1(sig_in[11]), .ip2(n22115), .ip3(n22114), 
        .ip4(n22113), .op(n22116) );
  or2_1 U26265 ( .ip1(n22117), .ip2(n22116), .op(n22118) );
  nand2_1 U26266 ( .ip1(n22123), .ip2(n22118), .op(n22170) );
  nand2_1 U26267 ( .ip1(n23938), .ip2(\x[111][14] ), .op(n22121) );
  nand2_1 U26268 ( .ip1(\x[111][12] ), .ip2(n24450), .op(n22120) );
  nand2_1 U26269 ( .ip1(\x[111][13] ), .ip2(n24235), .op(n22119) );
  nand3_1 U26270 ( .ip1(n22121), .ip2(n22120), .ip3(n22119), .op(n22122) );
  nand2_1 U26271 ( .ip1(n22123), .ip2(n22122), .op(n22216) );
  nand2_1 U26272 ( .ip1(n22170), .ip2(n22216), .op(n22124) );
  or2_1 U26273 ( .ip1(n22124), .ip2(n22174), .op(n22125) );
  nand2_1 U26274 ( .ip1(n22126), .ip2(n22125), .op(n22168) );
  inv_1 U26275 ( .ip(\x[110][11] ), .op(n22160) );
  and2_1 U26276 ( .ip1(n24451), .ip2(\x[110][10] ), .op(n22157) );
  inv_1 U26277 ( .ip(\x[110][9] ), .op(n22155) );
  and2_1 U26278 ( .ip1(n23804), .ip2(\x[110][8] ), .op(n22152) );
  inv_1 U26279 ( .ip(\x[110][5] ), .op(n22143) );
  nor2_1 U26280 ( .ip1(n22833), .ip2(n22143), .op(n22140) );
  inv_1 U26281 ( .ip(\x[110][3] ), .op(n22138) );
  inv_1 U26282 ( .ip(\x[110][1] ), .op(n22128) );
  nor2_1 U26283 ( .ip1(sig_in[1]), .ip2(n22128), .op(n22130) );
  inv_1 U26284 ( .ip(\x[110][0] ), .op(n22127) );
  not_ab_or_c_or_d U26285 ( .ip1(n24467), .ip2(n22128), .ip3(n23195), .ip4(
        n22127), .op(n22129) );
  not_ab_or_c_or_d U26286 ( .ip1(\x[110][2] ), .ip2(n24470), .ip3(n22130), 
        .ip4(n22129), .op(n22132) );
  nor2_1 U26287 ( .ip1(\x[110][2] ), .ip2(n24107), .op(n22131) );
  nor2_1 U26288 ( .ip1(n22132), .ip2(n22131), .op(n22133) );
  or2_1 U26289 ( .ip1(\x[110][3] ), .ip2(n22133), .op(n22135) );
  or2_1 U26290 ( .ip1(n24342), .ip2(n22133), .op(n22134) );
  nand2_1 U26291 ( .ip1(n22135), .ip2(n22134), .op(n22137) );
  nor2_1 U26292 ( .ip1(\x[110][4] ), .ip2(n24347), .op(n22136) );
  not_ab_or_c_or_d U26293 ( .ip1(n23251), .ip2(n22138), .ip3(n22137), .ip4(
        n22136), .op(n22139) );
  not_ab_or_c_or_d U26294 ( .ip1(\x[110][4] ), .ip2(n24347), .ip3(n22140), 
        .ip4(n22139), .op(n22142) );
  nor2_1 U26295 ( .ip1(\x[110][6] ), .ip2(n24355), .op(n22141) );
  not_ab_or_c_or_d U26296 ( .ip1(sig_in[5]), .ip2(n22143), .ip3(n22142), .ip4(
        n22141), .op(n22144) );
  or2_1 U26297 ( .ip1(\x[110][6] ), .ip2(n22144), .op(n22146) );
  or2_1 U26298 ( .ip1(n24485), .ip2(n22144), .op(n22145) );
  nand2_1 U26299 ( .ip1(n22146), .ip2(n22145), .op(n22147) );
  or2_1 U26300 ( .ip1(sig_in[7]), .ip2(n22147), .op(n22150) );
  inv_1 U26301 ( .ip(\x[110][7] ), .op(n22148) );
  or2_1 U26302 ( .ip1(n22148), .ip2(n22147), .op(n22149) );
  nand2_1 U26303 ( .ip1(n22150), .ip2(n22149), .op(n22151) );
  not_ab_or_c_or_d U26304 ( .ip1(\x[110][7] ), .ip2(n24142), .ip3(n22152), 
        .ip4(n22151), .op(n22154) );
  nor2_1 U26305 ( .ip1(\x[110][8] ), .ip2(n24100), .op(n22153) );
  not_ab_or_c_or_d U26306 ( .ip1(sig_in[9]), .ip2(n22155), .ip3(n22154), .ip4(
        n22153), .op(n22156) );
  not_ab_or_c_or_d U26307 ( .ip1(\x[110][9] ), .ip2(n24455), .ip3(n22157), 
        .ip4(n22156), .op(n22159) );
  nor2_1 U26308 ( .ip1(\x[110][10] ), .ip2(n24457), .op(n22158) );
  not_ab_or_c_or_d U26309 ( .ip1(sig_in[11]), .ip2(n22160), .ip3(n22159), 
        .ip4(n22158), .op(n22161) );
  or2_1 U26310 ( .ip1(\x[110][11] ), .ip2(n22161), .op(n22163) );
  or2_1 U26311 ( .ip1(n24371), .ip2(n22161), .op(n22162) );
  nand2_1 U26312 ( .ip1(n22163), .ip2(n22162), .op(n22279) );
  nor2_1 U26313 ( .ip1(\x[110][13] ), .ip2(n24137), .op(n22165) );
  nor2_1 U26314 ( .ip1(\x[110][12] ), .ip2(n24449), .op(n22164) );
  or2_1 U26315 ( .ip1(n22165), .ip2(n22164), .op(n22273) );
  or2_1 U26316 ( .ip1(n24185), .ip2(\x[110][14] ), .op(n22166) );
  nand2_1 U26317 ( .ip1(n22169), .ip2(n22166), .op(n22274) );
  nor3_1 U26318 ( .ip1(n22279), .ip2(n22273), .ip3(n22274), .op(n22167) );
  not_ab_or_c_or_d U26319 ( .ip1(n22169), .ip2(n22271), .ip3(n22168), .ip4(
        n22167), .op(n24592) );
  inv_1 U26320 ( .ip(n22170), .op(n22175) );
  nor2_1 U26321 ( .ip1(\x[112][15] ), .ip2(n24090), .op(n22177) );
  nor2_1 U26322 ( .ip1(\x[112][14] ), .ip2(n23938), .op(n22171) );
  or2_1 U26323 ( .ip1(\x[112][15] ), .ip2(n22171), .op(n22173) );
  or2_1 U26324 ( .ip1(n24384), .ip2(n22171), .op(n22172) );
  nand2_1 U26325 ( .ip1(n22173), .ip2(n22172), .op(n22267) );
  nor2_1 U26326 ( .ip1(n22177), .ip2(n22267), .op(n22260) );
  not_ab_or_c_or_d U26327 ( .ip1(n22176), .ip2(n22175), .ip3(n22260), .ip4(
        n22174), .op(n22218) );
  nand2_1 U26328 ( .ip1(n24327), .ip2(\x[112][14] ), .op(n22180) );
  inv_1 U26329 ( .ip(n22177), .op(n22179) );
  nand2_1 U26330 ( .ip1(\x[112][13] ), .ip2(n24235), .op(n22178) );
  nand3_1 U26331 ( .ip1(n22180), .ip2(n22179), .ip3(n22178), .op(n22214) );
  or2_1 U26332 ( .ip1(\x[112][12] ), .ip2(n22214), .op(n22182) );
  or2_1 U26333 ( .ip1(n24079), .ip2(n22214), .op(n22181) );
  nand2_1 U26334 ( .ip1(n22182), .ip2(n22181), .op(n22261) );
  nor2_1 U26335 ( .ip1(n21793), .ip2(\x[112][11] ), .op(n22210) );
  inv_1 U26336 ( .ip(\x[112][9] ), .op(n22206) );
  and2_1 U26337 ( .ip1(n23804), .ip2(\x[112][8] ), .op(n22203) );
  inv_1 U26338 ( .ip(\x[112][7] ), .op(n22201) );
  nor2_1 U26339 ( .ip1(n17732), .ip2(n22201), .op(n22198) );
  inv_1 U26340 ( .ip(\x[112][5] ), .op(n22196) );
  nor2_1 U26341 ( .ip1(sig_in[5]), .ip2(n22196), .op(n22193) );
  inv_1 U26342 ( .ip(\x[112][3] ), .op(n22191) );
  and2_1 U26343 ( .ip1(n24335), .ip2(\x[112][2] ), .op(n22188) );
  nand2_1 U26344 ( .ip1(\x[112][1] ), .ip2(n20652), .op(n22186) );
  nand2_1 U26345 ( .ip1(\x[112][0] ), .ip2(n24143), .op(n22185) );
  nor2_1 U26346 ( .ip1(\x[112][2] ), .ip2(n23659), .op(n22184) );
  nor2_1 U26347 ( .ip1(\x[112][1] ), .ip2(n20652), .op(n22183) );
  not_ab_or_c_or_d U26348 ( .ip1(n22186), .ip2(n22185), .ip3(n22184), .ip4(
        n22183), .op(n22187) );
  not_ab_or_c_or_d U26349 ( .ip1(\x[112][3] ), .ip2(n24342), .ip3(n22188), 
        .ip4(n22187), .op(n22190) );
  nor2_1 U26350 ( .ip1(\x[112][4] ), .ip2(n23721), .op(n22189) );
  not_ab_or_c_or_d U26351 ( .ip1(n23251), .ip2(n22191), .ip3(n22190), .ip4(
        n22189), .op(n22192) );
  not_ab_or_c_or_d U26352 ( .ip1(\x[112][4] ), .ip2(n24347), .ip3(n22193), 
        .ip4(n22192), .op(n22195) );
  nor2_1 U26353 ( .ip1(\x[112][6] ), .ip2(n24485), .op(n22194) );
  not_ab_or_c_or_d U26354 ( .ip1(sig_in[5]), .ip2(n22196), .ip3(n22195), .ip4(
        n22194), .op(n22197) );
  not_ab_or_c_or_d U26355 ( .ip1(\x[112][6] ), .ip2(n24355), .ip3(n22198), 
        .ip4(n22197), .op(n22200) );
  nor2_1 U26356 ( .ip1(\x[112][8] ), .ip2(n24358), .op(n22199) );
  not_ab_or_c_or_d U26357 ( .ip1(sig_in[7]), .ip2(n22201), .ip3(n22200), .ip4(
        n22199), .op(n22202) );
  not_ab_or_c_or_d U26358 ( .ip1(\x[112][9] ), .ip2(n24455), .ip3(n22203), 
        .ip4(n22202), .op(n22205) );
  nor2_1 U26359 ( .ip1(\x[112][10] ), .ip2(n23980), .op(n22204) );
  not_ab_or_c_or_d U26360 ( .ip1(sig_in[9]), .ip2(n22206), .ip3(n22205), .ip4(
        n22204), .op(n22208) );
  and2_1 U26361 ( .ip1(n24451), .ip2(\x[112][10] ), .op(n22207) );
  not_ab_or_c_or_d U26362 ( .ip1(\x[112][11] ), .ip2(n21793), .ip3(n22208), 
        .ip4(n22207), .op(n22209) );
  nor2_1 U26363 ( .ip1(n22210), .ip2(n22209), .op(n22265) );
  inv_1 U26364 ( .ip(n22265), .op(n22211) );
  nand2_1 U26365 ( .ip1(n22261), .ip2(n22211), .op(n22217) );
  nor2_1 U26366 ( .ip1(\x[112][13] ), .ip2(n24376), .op(n22213) );
  nor2_1 U26367 ( .ip1(\x[112][12] ), .ip2(n24450), .op(n22212) );
  nor2_1 U26368 ( .ip1(n22213), .ip2(n22212), .op(n22266) );
  or2_1 U26369 ( .ip1(n22214), .ip2(n22266), .op(n22215) );
  nand4_1 U26370 ( .ip1(n22218), .ip2(n22217), .ip3(n22216), .ip4(n22215), 
        .op(n26151) );
  nor2_1 U26371 ( .ip1(\x[113][9] ), .ip2(n24043), .op(n22239) );
  inv_1 U26372 ( .ip(\x[113][8] ), .op(n22219) );
  nor3_1 U26373 ( .ip1(sig_in[8]), .ip2(n22239), .ip3(n22219), .op(n22242) );
  and2_1 U26374 ( .ip1(n24461), .ip2(\x[113][7] ), .op(n22236) );
  inv_1 U26375 ( .ip(\x[113][5] ), .op(n22234) );
  nor2_1 U26376 ( .ip1(sig_in[5]), .ip2(n22234), .op(n22231) );
  nor2_1 U26377 ( .ip1(\x[113][4] ), .ip2(n24256), .op(n22229) );
  not_ab_or_c_or_d U26378 ( .ip1(\x[113][3] ), .ip2(n24476), .ip3(\x[113][2] ), 
        .ip4(n24470), .op(n22228) );
  nor2_1 U26379 ( .ip1(\x[113][3] ), .ip2(n24342), .op(n22227) );
  inv_1 U26380 ( .ip(\x[113][1] ), .op(n22221) );
  inv_1 U26381 ( .ip(\x[113][0] ), .op(n22220) );
  not_ab_or_c_or_d U26382 ( .ip1(n24467), .ip2(n22221), .ip3(n23195), .ip4(
        n22220), .op(n22225) );
  nand2_1 U26383 ( .ip1(\x[113][3] ), .ip2(n24476), .op(n22223) );
  nand2_1 U26384 ( .ip1(\x[113][1] ), .ip2(n21685), .op(n22222) );
  nand2_1 U26385 ( .ip1(n22223), .ip2(n22222), .op(n22224) );
  not_ab_or_c_or_d U26386 ( .ip1(\x[113][2] ), .ip2(n24470), .ip3(n22225), 
        .ip4(n22224), .op(n22226) );
  nor4_1 U26387 ( .ip1(n22229), .ip2(n22228), .ip3(n22227), .ip4(n22226), .op(
        n22230) );
  not_ab_or_c_or_d U26388 ( .ip1(\x[113][4] ), .ip2(n23860), .ip3(n22231), 
        .ip4(n22230), .op(n22233) );
  nor2_1 U26389 ( .ip1(\x[113][6] ), .ip2(n23509), .op(n22232) );
  not_ab_or_c_or_d U26390 ( .ip1(sig_in[5]), .ip2(n22234), .ip3(n22233), .ip4(
        n22232), .op(n22235) );
  not_ab_or_c_or_d U26391 ( .ip1(\x[113][6] ), .ip2(n24045), .ip3(n22236), 
        .ip4(n22235), .op(n22240) );
  nor2_1 U26392 ( .ip1(\x[113][7] ), .ip2(n24044), .op(n22238) );
  nor2_1 U26393 ( .ip1(\x[113][8] ), .ip2(n24358), .op(n22237) );
  nor4_1 U26394 ( .ip1(n22240), .ip2(n22239), .ip3(n22238), .ip4(n22237), .op(
        n22241) );
  not_ab_or_c_or_d U26395 ( .ip1(\x[113][10] ), .ip2(n24370), .ip3(n22242), 
        .ip4(n22241), .op(n22246) );
  nand2_1 U26396 ( .ip1(\x[113][9] ), .ip2(n24043), .op(n22245) );
  nor2_1 U26397 ( .ip1(\x[113][10] ), .ip2(n23980), .op(n22244) );
  nor2_1 U26398 ( .ip1(\x[113][11] ), .ip2(n24371), .op(n22243) );
  not_ab_or_c_or_d U26399 ( .ip1(n22246), .ip2(n22245), .ip3(n22244), .ip4(
        n22243), .op(n22247) );
  or2_1 U26400 ( .ip1(\x[113][11] ), .ip2(n22247), .op(n22249) );
  or2_1 U26401 ( .ip1(n24239), .ip2(n22247), .op(n22248) );
  nand2_1 U26402 ( .ip1(n22249), .ip2(n22248), .op(n22784) );
  and2_1 U26403 ( .ip1(n23895), .ip2(\x[113][13] ), .op(n22250) );
  nor2_1 U26404 ( .ip1(\x[113][15] ), .ip2(n24090), .op(n22259) );
  not_ab_or_c_or_d U26405 ( .ip1(\x[113][14] ), .ip2(n24327), .ip3(n22250), 
        .ip4(n22259), .op(n22264) );
  inv_1 U26406 ( .ip(n22264), .op(n22251) );
  or2_1 U26407 ( .ip1(\x[113][12] ), .ip2(n22251), .op(n22253) );
  or2_1 U26408 ( .ip1(n24449), .ip2(n22251), .op(n22252) );
  nand2_1 U26409 ( .ip1(n22253), .ip2(n22252), .op(n22778) );
  nand2_1 U26410 ( .ip1(n22784), .ip2(n22778), .op(n22270) );
  nor2_1 U26411 ( .ip1(\x[113][13] ), .ip2(n24137), .op(n22255) );
  nor2_1 U26412 ( .ip1(\x[113][12] ), .ip2(n24079), .op(n22254) );
  or2_1 U26413 ( .ip1(n22255), .ip2(n22254), .op(n22782) );
  and2_1 U26414 ( .ip1(n24186), .ip2(\x[113][15] ), .op(n22779) );
  or2_1 U26415 ( .ip1(sig_in[14]), .ip2(n22779), .op(n22258) );
  inv_1 U26416 ( .ip(\x[113][14] ), .op(n22256) );
  or2_1 U26417 ( .ip1(n22256), .ip2(n22779), .op(n22257) );
  nand2_1 U26418 ( .ip1(n22258), .ip2(n22257), .op(n22781) );
  nor2_1 U26419 ( .ip1(n22259), .ip2(n22781), .op(n22263) );
  nor2_1 U26420 ( .ip1(n22261), .ip2(n22260), .op(n22262) );
  not_ab_or_c_or_d U26421 ( .ip1(n22264), .ip2(n22782), .ip3(n22263), .ip4(
        n22262), .op(n22269) );
  nand3_1 U26422 ( .ip1(n22267), .ip2(n22266), .ip3(n22265), .op(n22268) );
  nand3_1 U26423 ( .ip1(n22270), .ip2(n22269), .ip3(n22268), .op(n26152) );
  nand2_1 U26424 ( .ip1(n26151), .ip2(n26152), .op(n24594) );
  nor2_1 U26425 ( .ip1(n24592), .ip2(n24594), .op(n24595) );
  inv_1 U26426 ( .ip(n22271), .op(n22280) );
  and2_1 U26427 ( .ip1(n22273), .ip2(n22272), .op(n22278) );
  inv_1 U26428 ( .ip(n22274), .op(n22276) );
  nor2_1 U26429 ( .ip1(n22276), .ip2(n22275), .op(n22277) );
  not_ab_or_c_or_d U26430 ( .ip1(n22280), .ip2(n22279), .ip3(n22278), .ip4(
        n22277), .op(n22291) );
  nand3_1 U26431 ( .ip1(n22284), .ip2(n22282), .ip3(n22281), .op(n22290) );
  nand2_1 U26432 ( .ip1(n22284), .ip2(n22283), .op(n22289) );
  inv_1 U26433 ( .ip(n22285), .op(n22286) );
  nand2_1 U26434 ( .ip1(n22287), .ip2(n22286), .op(n22288) );
  nand4_1 U26435 ( .ip1(n22291), .ip2(n22290), .ip3(n22289), .ip4(n22288), 
        .op(n24596) );
  nand2_1 U26436 ( .ip1(n24595), .ip2(n24596), .op(n24959) );
  nor2_1 U26437 ( .ip1(n24960), .ip2(n24959), .op(n24586) );
  inv_1 U26438 ( .ip(n22292), .op(n22296) );
  or2_1 U26439 ( .ip1(n22293), .ip2(n22296), .op(n22299) );
  nand2_1 U26440 ( .ip1(n22295), .ip2(n22294), .op(n22297) );
  or2_1 U26441 ( .ip1(n22297), .ip2(n22296), .op(n22298) );
  nand2_1 U26442 ( .ip1(n22299), .ip2(n22298), .op(n22307) );
  inv_1 U26443 ( .ip(n22300), .op(n22302) );
  nor2_1 U26444 ( .ip1(n22302), .ip2(n22301), .op(n22306) );
  and2_1 U26445 ( .ip1(n22304), .ip2(n22303), .op(n22305) );
  or4_1 U26446 ( .ip1(n22308), .ip2(n22307), .ip3(n22306), .ip4(n22305), .op(
        n24587) );
  nand2_1 U26447 ( .ip1(n24586), .ip2(n24587), .op(n24522) );
  nor2_1 U26448 ( .ip1(n24524), .ip2(n24522), .op(n24583) );
  inv_1 U26449 ( .ip(n22319), .op(n22310) );
  nand2_1 U26450 ( .ip1(n22310), .ip2(n22309), .op(n22347) );
  inv_1 U26451 ( .ip(n22311), .op(n22313) );
  nand2_1 U26452 ( .ip1(\x[106][8] ), .ip2(n23971), .op(n22312) );
  nand2_1 U26453 ( .ip1(n22313), .ip2(n22312), .op(n22315) );
  nand2_1 U26454 ( .ip1(n22315), .ip2(n22314), .op(n22317) );
  nand2_1 U26455 ( .ip1(n22317), .ip2(n22316), .op(n22320) );
  not_ab_or_c_or_d U26456 ( .ip1(n22321), .ip2(n22320), .ip3(n22319), .ip4(
        n22318), .op(n22342) );
  or3_1 U26457 ( .ip1(n23779), .ip2(n22323), .ip3(n22322), .op(n22324) );
  nand2_1 U26458 ( .ip1(n22325), .ip2(n22324), .op(n22326) );
  nand2_1 U26459 ( .ip1(n22327), .ip2(n22326), .op(n22336) );
  inv_1 U26460 ( .ip(n22328), .op(n22329) );
  nand3_1 U26461 ( .ip1(n22331), .ip2(n22330), .ip3(n22329), .op(n22335) );
  nor2_1 U26462 ( .ip1(\x[105][14] ), .ip2(n23938), .op(n22334) );
  inv_1 U26463 ( .ip(n22332), .op(n22333) );
  not_ab_or_c_or_d U26464 ( .ip1(n22336), .ip2(n22335), .ip3(n22334), .ip4(
        n22333), .op(n22338) );
  not_ab_or_c_or_d U26465 ( .ip1(\x[105][14] ), .ip2(n24230), .ip3(n22338), 
        .ip4(n22337), .op(n22339) );
  nor2_1 U26466 ( .ip1(n22340), .ip2(n22339), .op(n22341) );
  not_ab_or_c_or_d U26467 ( .ip1(n22344), .ip2(n22343), .ip3(n22342), .ip4(
        n22341), .op(n22346) );
  nand3_1 U26468 ( .ip1(n22347), .ip2(n22346), .ip3(n22345), .op(n24584) );
  nand2_1 U26469 ( .ip1(n24583), .ip2(n24584), .op(n24590) );
  nor2_1 U26470 ( .ip1(n24589), .ip2(n24590), .op(n24610) );
  inv_1 U26471 ( .ip(n22348), .op(n22349) );
  nand2_1 U26472 ( .ip1(n22350), .ip2(n22349), .op(n22366) );
  nand2_1 U26473 ( .ip1(n22352), .ip2(n22351), .op(n22354) );
  nand2_1 U26474 ( .ip1(n22354), .ip2(n22353), .op(n22356) );
  nand2_1 U26475 ( .ip1(n22356), .ip2(n22355), .op(n22365) );
  inv_1 U26476 ( .ip(n22357), .op(n22361) );
  nand2_1 U26477 ( .ip1(n22359), .ip2(n22358), .op(n22360) );
  nand2_1 U26478 ( .ip1(n22361), .ip2(n22360), .op(n22362) );
  nand2_1 U26479 ( .ip1(n22363), .ip2(n22362), .op(n22364) );
  nand3_1 U26480 ( .ip1(n22366), .ip2(n22365), .ip3(n22364), .op(n24612) );
  nand2_1 U26481 ( .ip1(n24610), .ip2(n24612), .op(n24582) );
  nor2_1 U26482 ( .ip1(n24580), .ip2(n24582), .op(n24607) );
  inv_1 U26483 ( .ip(n22367), .op(n22369) );
  nand2_1 U26484 ( .ip1(n22369), .ip2(n22368), .op(n22383) );
  inv_1 U26485 ( .ip(n22370), .op(n22376) );
  inv_1 U26486 ( .ip(n22371), .op(n22375) );
  nor2_1 U26487 ( .ip1(n22373), .ip2(n22372), .op(n22374) );
  not_ab_or_c_or_d U26488 ( .ip1(n22377), .ip2(n22376), .ip3(n22375), .ip4(
        n22374), .op(n22382) );
  nand3_1 U26489 ( .ip1(n22380), .ip2(n22379), .ip3(n22378), .op(n22381) );
  nand3_1 U26490 ( .ip1(n22383), .ip2(n22382), .ip3(n22381), .op(n24608) );
  nand2_1 U26491 ( .ip1(n24607), .ip2(n24608), .op(n24606) );
  nor2_1 U26492 ( .ip1(n24604), .ip2(n24606), .op(n24525) );
  inv_1 U26493 ( .ip(n22384), .op(n22399) );
  inv_1 U26494 ( .ip(n22385), .op(n22398) );
  inv_1 U26495 ( .ip(n22386), .op(n22389) );
  inv_1 U26496 ( .ip(n22387), .op(n22388) );
  not_ab_or_c_or_d U26497 ( .ip1(n22391), .ip2(n22390), .ip3(n22389), .ip4(
        n22388), .op(n22392) );
  nor2_1 U26498 ( .ip1(n22393), .ip2(n22392), .op(n22396) );
  nand2_1 U26499 ( .ip1(n22399), .ip2(n22394), .op(n22395) );
  nor2_1 U26500 ( .ip1(n22396), .ip2(n22395), .op(n22397) );
  ab_or_c_or_d U26501 ( .ip1(n22400), .ip2(n22399), .ip3(n22398), .ip4(n22397), 
        .op(n27367) );
  nand2_1 U26502 ( .ip1(n24525), .ip2(n27367), .op(n27142) );
  and2_1 U26503 ( .ip1(n24332), .ip2(\x[114][13] ), .op(n22401) );
  nor2_1 U26504 ( .ip1(\x[114][15] ), .ip2(n24090), .op(n22406) );
  not_ab_or_c_or_d U26505 ( .ip1(\x[114][14] ), .ip2(n24230), .ip3(n22401), 
        .ip4(n22406), .op(n22788) );
  nand2_1 U26506 ( .ip1(\x[114][12] ), .ip2(n24449), .op(n22402) );
  nand2_1 U26507 ( .ip1(n22788), .ip2(n22402), .op(n22790) );
  nor2_1 U26508 ( .ip1(\x[114][14] ), .ip2(n24230), .op(n22403) );
  or2_1 U26509 ( .ip1(\x[114][15] ), .ip2(n22403), .op(n22405) );
  or2_1 U26510 ( .ip1(n24384), .ip2(n22403), .op(n22404) );
  nand2_1 U26511 ( .ip1(n22405), .ip2(n22404), .op(n22445) );
  nor2_1 U26512 ( .ip1(n22406), .ip2(n22445), .op(n22785) );
  inv_1 U26513 ( .ip(n22785), .op(n22498) );
  nor2_1 U26514 ( .ip1(\x[114][13] ), .ip2(n24137), .op(n22407) );
  or2_1 U26515 ( .ip1(n17845), .ip2(n22407), .op(n22410) );
  inv_1 U26516 ( .ip(\x[114][12] ), .op(n22408) );
  or2_1 U26517 ( .ip1(n22408), .ip2(n22407), .op(n22409) );
  nand2_1 U26518 ( .ip1(n22410), .ip2(n22409), .op(n22780) );
  inv_1 U26519 ( .ip(\x[114][7] ), .op(n22428) );
  nor2_1 U26520 ( .ip1(n22428), .ip2(n17732), .op(n22430) );
  nor2_1 U26521 ( .ip1(\x[114][6] ), .ip2(n24355), .op(n22427) );
  and2_1 U26522 ( .ip1(n24107), .ip2(\x[114][2] ), .op(n22416) );
  nand2_1 U26523 ( .ip1(\x[114][1] ), .ip2(n20652), .op(n22414) );
  nand2_1 U26524 ( .ip1(\x[114][0] ), .ip2(n24143), .op(n22413) );
  nor2_1 U26525 ( .ip1(\x[114][2] ), .ip2(n23659), .op(n22412) );
  nor2_1 U26526 ( .ip1(\x[114][1] ), .ip2(n21685), .op(n22411) );
  not_ab_or_c_or_d U26527 ( .ip1(n22414), .ip2(n22413), .ip3(n22412), .ip4(
        n22411), .op(n22415) );
  not_ab_or_c_or_d U26528 ( .ip1(\x[114][3] ), .ip2(n24476), .ip3(n22416), 
        .ip4(n22415), .op(n22419) );
  nor2_1 U26529 ( .ip1(\x[114][5] ), .ip2(n24482), .op(n22420) );
  nor2_1 U26530 ( .ip1(\x[114][3] ), .ip2(n24342), .op(n22418) );
  nor2_1 U26531 ( .ip1(\x[114][4] ), .ip2(n23860), .op(n22417) );
  nor4_1 U26532 ( .ip1(n22419), .ip2(n22420), .ip3(n22418), .ip4(n22417), .op(
        n22425) );
  inv_1 U26533 ( .ip(n22420), .op(n22421) );
  nand3_1 U26534 ( .ip1(n23721), .ip2(\x[114][4] ), .ip3(n22421), .op(n22423)
         );
  nand2_1 U26535 ( .ip1(\x[114][6] ), .ip2(n24485), .op(n22422) );
  nand2_1 U26536 ( .ip1(n22423), .ip2(n22422), .op(n22424) );
  not_ab_or_c_or_d U26537 ( .ip1(\x[114][5] ), .ip2(n24482), .ip3(n22425), 
        .ip4(n22424), .op(n22426) );
  not_ab_or_c_or_d U26538 ( .ip1(sig_in[7]), .ip2(n22428), .ip3(n22427), .ip4(
        n22426), .op(n22429) );
  or2_1 U26539 ( .ip1(n22430), .ip2(n22429), .op(n22434) );
  nand2_1 U26540 ( .ip1(n22434), .ip2(\x[114][8] ), .op(n22437) );
  nor2_1 U26541 ( .ip1(\x[114][11] ), .ip2(n24456), .op(n22439) );
  or2_1 U26542 ( .ip1(sig_in[10]), .ip2(n22439), .op(n22432) );
  inv_1 U26543 ( .ip(\x[114][10] ), .op(n22440) );
  or2_1 U26544 ( .ip1(n22440), .ip2(n22439), .op(n22431) );
  nand2_1 U26545 ( .ip1(n22432), .ip2(n22431), .op(n22438) );
  or2_1 U26546 ( .ip1(n23981), .ip2(\x[114][9] ), .op(n22433) );
  nand2_1 U26547 ( .ip1(n22438), .ip2(n22433), .op(n22436) );
  nor2_1 U26548 ( .ip1(n22434), .ip2(\x[114][8] ), .op(n22435) );
  ab_or_c_or_d U26549 ( .ip1(n23779), .ip2(n22437), .ip3(n22436), .ip4(n22435), 
        .op(n22444) );
  nand3_1 U26550 ( .ip1(\x[114][9] ), .ip2(n22438), .ip3(n24269), .op(n22443)
         );
  nand2_1 U26551 ( .ip1(\x[114][11] ), .ip2(n24239), .op(n22442) );
  or3_1 U26552 ( .ip1(n22440), .ip2(sig_in[10]), .ip3(n22439), .op(n22441) );
  nand4_1 U26553 ( .ip1(n22444), .ip2(n22443), .ip3(n22442), .ip4(n22441), 
        .op(n22789) );
  and3_1 U26554 ( .ip1(n22780), .ip2(n22445), .ip3(n22789), .op(n22497) );
  nor2_1 U26555 ( .ip1(\x[115][13] ), .ip2(n24137), .op(n22446) );
  or2_1 U26556 ( .ip1(sig_in[12]), .ip2(n22446), .op(n22449) );
  inv_1 U26557 ( .ip(\x[115][12] ), .op(n22447) );
  or2_1 U26558 ( .ip1(n22447), .ip2(n22446), .op(n22448) );
  nand2_1 U26559 ( .ip1(n22449), .ip2(n22448), .op(n22773) );
  nor2_1 U26560 ( .ip1(\x[115][15] ), .ip2(n24090), .op(n22774) );
  or2_1 U26561 ( .ip1(n22773), .ip2(n22774), .op(n22495) );
  inv_1 U26562 ( .ip(\x[115][11] ), .op(n22485) );
  and2_1 U26563 ( .ip1(n24451), .ip2(\x[115][10] ), .op(n22481) );
  inv_1 U26564 ( .ip(\x[115][9] ), .op(n22479) );
  and2_1 U26565 ( .ip1(n24491), .ip2(\x[115][8] ), .op(n22471) );
  inv_1 U26566 ( .ip(\x[115][6] ), .op(n22469) );
  nor2_1 U26567 ( .ip1(\x[115][5] ), .ip2(n24350), .op(n22463) );
  and2_1 U26568 ( .ip1(n24347), .ip2(\x[115][4] ), .op(n22461) );
  inv_1 U26569 ( .ip(\x[115][3] ), .op(n22458) );
  and2_1 U26570 ( .ip1(n24335), .ip2(\x[115][2] ), .op(n22455) );
  nand2_1 U26571 ( .ip1(\x[115][1] ), .ip2(n21685), .op(n22453) );
  nand2_1 U26572 ( .ip1(\x[115][0] ), .ip2(n24143), .op(n22452) );
  nor2_1 U26573 ( .ip1(\x[115][2] ), .ip2(n23659), .op(n22451) );
  nor2_1 U26574 ( .ip1(\x[115][1] ), .ip2(n20652), .op(n22450) );
  not_ab_or_c_or_d U26575 ( .ip1(n22453), .ip2(n22452), .ip3(n22451), .ip4(
        n22450), .op(n22454) );
  not_ab_or_c_or_d U26576 ( .ip1(\x[115][3] ), .ip2(n24342), .ip3(n22455), 
        .ip4(n22454), .op(n22457) );
  nor2_1 U26577 ( .ip1(\x[115][4] ), .ip2(n24347), .op(n22456) );
  not_ab_or_c_or_d U26578 ( .ip1(n23251), .ip2(n22458), .ip3(n22457), .ip4(
        n22456), .op(n22460) );
  and2_1 U26579 ( .ip1(n24119), .ip2(\x[115][5] ), .op(n22459) );
  nor3_1 U26580 ( .ip1(n22461), .ip2(n22460), .ip3(n22459), .op(n22462) );
  nor2_1 U26581 ( .ip1(n22463), .ip2(n22462), .op(n22464) );
  or2_1 U26582 ( .ip1(\x[115][6] ), .ip2(n22464), .op(n22466) );
  or2_1 U26583 ( .ip1(n24355), .ip2(n22464), .op(n22465) );
  nand2_1 U26584 ( .ip1(n22466), .ip2(n22465), .op(n22468) );
  nor2_1 U26585 ( .ip1(\x[115][7] ), .ip2(n24044), .op(n22467) );
  not_ab_or_c_or_d U26586 ( .ip1(sig_in[6]), .ip2(n22469), .ip3(n22468), .ip4(
        n22467), .op(n22470) );
  not_ab_or_c_or_d U26587 ( .ip1(\x[115][7] ), .ip2(n24142), .ip3(n22471), 
        .ip4(n22470), .op(n22473) );
  nor2_1 U26588 ( .ip1(\x[115][8] ), .ip2(n23971), .op(n22472) );
  nor2_1 U26589 ( .ip1(n22473), .ip2(n22472), .op(n22474) );
  or2_1 U26590 ( .ip1(\x[115][9] ), .ip2(n22474), .op(n22476) );
  or2_1 U26591 ( .ip1(n24455), .ip2(n22474), .op(n22475) );
  nand2_1 U26592 ( .ip1(n22476), .ip2(n22475), .op(n22478) );
  nor2_1 U26593 ( .ip1(\x[115][10] ), .ip2(n23980), .op(n22477) );
  not_ab_or_c_or_d U26594 ( .ip1(sig_in[9]), .ip2(n22479), .ip3(n22478), .ip4(
        n22477), .op(n22480) );
  not_ab_or_c_or_d U26595 ( .ip1(\x[115][11] ), .ip2(n24456), .ip3(n22481), 
        .ip4(n22480), .op(n22484) );
  or2_1 U26596 ( .ip1(n24185), .ip2(\x[115][14] ), .op(n22483) );
  nand2_1 U26597 ( .ip1(\x[115][15] ), .ip2(n24329), .op(n22482) );
  nand2_1 U26598 ( .ip1(n22483), .ip2(n22482), .op(n22486) );
  not_ab_or_c_or_d U26599 ( .ip1(sig_in[11]), .ip2(n22485), .ip3(n22484), 
        .ip4(n22486), .op(n22772) );
  inv_1 U26600 ( .ip(n22772), .op(n22492) );
  inv_1 U26601 ( .ip(n22486), .op(n22491) );
  nand2_1 U26602 ( .ip1(n24230), .ip2(\x[115][14] ), .op(n22489) );
  nand2_1 U26603 ( .ip1(\x[115][12] ), .ip2(n24450), .op(n22488) );
  nand2_1 U26604 ( .ip1(\x[115][13] ), .ip2(n24081), .op(n22487) );
  nand3_1 U26605 ( .ip1(n22489), .ip2(n22488), .ip3(n22487), .op(n22490) );
  nand2_1 U26606 ( .ip1(n22491), .ip2(n22490), .op(n22775) );
  nand2_1 U26607 ( .ip1(n22492), .ip2(n22775), .op(n22493) );
  or2_1 U26608 ( .ip1(n22493), .ip2(n22774), .op(n22494) );
  nand2_1 U26609 ( .ip1(n22495), .ip2(n22494), .op(n22496) );
  not_ab_or_c_or_d U26610 ( .ip1(n22790), .ip2(n22498), .ip3(n22497), .ip4(
        n22496), .op(n24639) );
  nand2_1 U26611 ( .ip1(n24384), .ip2(\x[117][15] ), .op(n22752) );
  inv_1 U26612 ( .ip(n22752), .op(n22499) );
  or2_1 U26613 ( .ip1(sig_in[14]), .ip2(n22499), .op(n22502) );
  inv_1 U26614 ( .ip(\x[117][14] ), .op(n22500) );
  or2_1 U26615 ( .ip1(n22500), .ip2(n22499), .op(n22501) );
  nand2_1 U26616 ( .ip1(n22502), .ip2(n22501), .op(n22740) );
  nor2_1 U26617 ( .ip1(\x[117][15] ), .ip2(n24090), .op(n22589) );
  nor2_1 U26618 ( .ip1(n22740), .ip2(n22589), .op(n22597) );
  nand2_1 U26619 ( .ip1(n24382), .ip2(\x[116][14] ), .op(n22505) );
  nor2_1 U26620 ( .ip1(n24384), .ip2(\x[116][15] ), .op(n22511) );
  inv_1 U26621 ( .ip(n22511), .op(n22504) );
  nand2_1 U26622 ( .ip1(\x[116][13] ), .ip2(n24235), .op(n22503) );
  nand3_1 U26623 ( .ip1(n22505), .ip2(n22504), .ip3(n22503), .op(n22765) );
  or2_1 U26624 ( .ip1(\x[116][12] ), .ip2(n22765), .op(n22507) );
  or2_1 U26625 ( .ip1(n24079), .ip2(n22765), .op(n22506) );
  nand2_1 U26626 ( .ip1(n22507), .ip2(n22506), .op(n22762) );
  nor2_1 U26627 ( .ip1(\x[116][14] ), .ip2(n24230), .op(n22508) );
  or2_1 U26628 ( .ip1(\x[116][15] ), .ip2(n22508), .op(n22510) );
  or2_1 U26629 ( .ip1(n24384), .ip2(n22508), .op(n22509) );
  nand2_1 U26630 ( .ip1(n22510), .ip2(n22509), .op(n22548) );
  nor2_1 U26631 ( .ip1(n22511), .ip2(n22548), .op(n22766) );
  nor2_1 U26632 ( .ip1(n22762), .ip2(n22766), .op(n22596) );
  nand2_1 U26633 ( .ip1(\x[116][10] ), .ip2(n23146), .op(n22539) );
  nor2_1 U26634 ( .ip1(\x[116][9] ), .ip2(n24043), .op(n22534) );
  inv_1 U26635 ( .ip(\x[116][8] ), .op(n22512) );
  nor3_1 U26636 ( .ip1(sig_in[8]), .ip2(n22534), .ip3(n22512), .op(n22537) );
  and2_1 U26637 ( .ip1(n24461), .ip2(\x[116][7] ), .op(n22531) );
  inv_1 U26638 ( .ip(\x[116][3] ), .op(n22520) );
  inv_1 U26639 ( .ip(\x[116][1] ), .op(n22515) );
  nor2_1 U26640 ( .ip1(n22513), .ip2(n22515), .op(n22517) );
  inv_1 U26641 ( .ip(\x[116][0] ), .op(n22514) );
  not_ab_or_c_or_d U26642 ( .ip1(n24467), .ip2(n22515), .ip3(n23195), .ip4(
        n22514), .op(n22516) );
  not_ab_or_c_or_d U26643 ( .ip1(\x[116][2] ), .ip2(n24470), .ip3(n22517), 
        .ip4(n22516), .op(n22519) );
  nor2_1 U26644 ( .ip1(\x[116][2] ), .ip2(n23659), .op(n22518) );
  not_ab_or_c_or_d U26645 ( .ip1(sig_in[3]), .ip2(n22520), .ip3(n22519), .ip4(
        n22518), .op(n22524) );
  nand2_1 U26646 ( .ip1(\x[116][5] ), .ip2(n24119), .op(n22522) );
  nand2_1 U26647 ( .ip1(\x[116][4] ), .ip2(n23721), .op(n22521) );
  nand2_1 U26648 ( .ip1(n22522), .ip2(n22521), .op(n22523) );
  not_ab_or_c_or_d U26649 ( .ip1(\x[116][3] ), .ip2(n22525), .ip3(n22524), 
        .ip4(n22523), .op(n22529) );
  nor2_1 U26650 ( .ip1(\x[116][6] ), .ip2(n23770), .op(n22528) );
  nor2_1 U26651 ( .ip1(\x[116][5] ), .ip2(n24350), .op(n22527) );
  not_ab_or_c_or_d U26652 ( .ip1(\x[116][5] ), .ip2(n23600), .ip3(\x[116][4] ), 
        .ip4(n24256), .op(n22526) );
  nor4_1 U26653 ( .ip1(n22529), .ip2(n22528), .ip3(n22527), .ip4(n22526), .op(
        n22530) );
  not_ab_or_c_or_d U26654 ( .ip1(\x[116][6] ), .ip2(n24045), .ip3(n22531), 
        .ip4(n22530), .op(n22535) );
  nor2_1 U26655 ( .ip1(\x[116][7] ), .ip2(n24044), .op(n22533) );
  nor2_1 U26656 ( .ip1(\x[116][8] ), .ip2(n24100), .op(n22532) );
  nor4_1 U26657 ( .ip1(n22535), .ip2(n22534), .ip3(n22533), .ip4(n22532), .op(
        n22536) );
  not_ab_or_c_or_d U26658 ( .ip1(\x[116][9] ), .ip2(n24455), .ip3(n22537), 
        .ip4(n22536), .op(n22538) );
  nand2_1 U26659 ( .ip1(n22539), .ip2(n22538), .op(n22545) );
  nor2_1 U26660 ( .ip1(\x[116][10] ), .ip2(n23980), .op(n22540) );
  or2_1 U26661 ( .ip1(sig_in[11]), .ip2(n22540), .op(n22543) );
  inv_1 U26662 ( .ip(\x[116][11] ), .op(n22541) );
  or2_1 U26663 ( .ip1(n22541), .ip2(n22540), .op(n22542) );
  nand2_1 U26664 ( .ip1(n22543), .ip2(n22542), .op(n22544) );
  nand2_1 U26665 ( .ip1(n22545), .ip2(n22544), .op(n22547) );
  nand2_1 U26666 ( .ip1(\x[116][11] ), .ip2(n24239), .op(n22546) );
  nand2_1 U26667 ( .ip1(n22547), .ip2(n22546), .op(n22764) );
  inv_1 U26668 ( .ip(\x[116][12] ), .op(n22551) );
  nor2_1 U26669 ( .ip1(\x[116][13] ), .ip2(n24081), .op(n22550) );
  inv_1 U26670 ( .ip(n22548), .op(n22549) );
  not_ab_or_c_or_d U26671 ( .ip1(sig_in[12]), .ip2(n22551), .ip3(n22550), 
        .ip4(n22549), .op(n22769) );
  and2_1 U26672 ( .ip1(n22764), .ip2(n22769), .op(n22595) );
  nor2_1 U26673 ( .ip1(\x[117][13] ), .ip2(n24137), .op(n22552) );
  or2_1 U26674 ( .ip1(sig_in[12]), .ip2(n22552), .op(n22555) );
  inv_1 U26675 ( .ip(\x[117][12] ), .op(n22553) );
  or2_1 U26676 ( .ip1(n22553), .ip2(n22552), .op(n22554) );
  nand2_1 U26677 ( .ip1(n22555), .ip2(n22554), .op(n22745) );
  nand2_1 U26678 ( .ip1(\x[117][9] ), .ip2(n24043), .op(n22558) );
  nor2_1 U26679 ( .ip1(\x[117][11] ), .ip2(n21793), .op(n22557) );
  nor2_1 U26680 ( .ip1(\x[117][10] ), .ip2(n23980), .op(n22556) );
  or2_1 U26681 ( .ip1(n22557), .ip2(n22556), .op(n22562) );
  or2_1 U26682 ( .ip1(n22558), .ip2(n22562), .op(n22561) );
  nand2_1 U26683 ( .ip1(\x[117][10] ), .ip2(n23146), .op(n22559) );
  or2_1 U26684 ( .ip1(n22559), .ip2(n22562), .op(n22560) );
  nand2_1 U26685 ( .ip1(n22561), .ip2(n22560), .op(n22588) );
  nor2_1 U26686 ( .ip1(n24455), .ip2(\x[117][9] ), .op(n22563) );
  nor2_1 U26687 ( .ip1(n22563), .ip2(n22562), .op(n22584) );
  inv_1 U26688 ( .ip(\x[117][7] ), .op(n22582) );
  nor2_1 U26689 ( .ip1(n17732), .ip2(n22582), .op(n22579) );
  inv_1 U26690 ( .ip(\x[117][5] ), .op(n22577) );
  nor2_1 U26691 ( .ip1(sig_in[5]), .ip2(n22577), .op(n22574) );
  inv_1 U26692 ( .ip(\x[117][3] ), .op(n22572) );
  and2_1 U26693 ( .ip1(n24107), .ip2(\x[117][2] ), .op(n22569) );
  nand2_1 U26694 ( .ip1(\x[117][1] ), .ip2(n20652), .op(n22567) );
  nand2_1 U26695 ( .ip1(\x[117][0] ), .ip2(n24143), .op(n22566) );
  nor2_1 U26696 ( .ip1(\x[117][2] ), .ip2(n23659), .op(n22565) );
  nor2_1 U26697 ( .ip1(\x[117][1] ), .ip2(n21685), .op(n22564) );
  not_ab_or_c_or_d U26698 ( .ip1(n22567), .ip2(n22566), .ip3(n22565), .ip4(
        n22564), .op(n22568) );
  not_ab_or_c_or_d U26699 ( .ip1(\x[117][3] ), .ip2(n24342), .ip3(n22569), 
        .ip4(n22568), .op(n22571) );
  nor2_1 U26700 ( .ip1(\x[117][4] ), .ip2(n23721), .op(n22570) );
  not_ab_or_c_or_d U26701 ( .ip1(sig_in[3]), .ip2(n22572), .ip3(n22571), .ip4(
        n22570), .op(n22573) );
  not_ab_or_c_or_d U26702 ( .ip1(\x[117][4] ), .ip2(n23860), .ip3(n22574), 
        .ip4(n22573), .op(n22576) );
  nor2_1 U26703 ( .ip1(\x[117][6] ), .ip2(n24485), .op(n22575) );
  not_ab_or_c_or_d U26704 ( .ip1(sig_in[5]), .ip2(n22577), .ip3(n22576), .ip4(
        n22575), .op(n22578) );
  not_ab_or_c_or_d U26705 ( .ip1(\x[117][6] ), .ip2(n24045), .ip3(n22579), 
        .ip4(n22578), .op(n22581) );
  nor2_1 U26706 ( .ip1(\x[117][8] ), .ip2(n23971), .op(n22580) );
  not_ab_or_c_or_d U26707 ( .ip1(sig_in[7]), .ip2(n22582), .ip3(n22581), .ip4(
        n22580), .op(n22583) );
  nand2_1 U26708 ( .ip1(n22584), .ip2(n22583), .op(n22586) );
  nand3_1 U26709 ( .ip1(n22584), .ip2(n23971), .ip3(\x[117][8] ), .op(n22585)
         );
  nand2_1 U26710 ( .ip1(n22586), .ip2(n22585), .op(n22587) );
  not_ab_or_c_or_d U26711 ( .ip1(\x[117][11] ), .ip2(n24136), .ip3(n22588), 
        .ip4(n22587), .op(n22748) );
  nand2_1 U26712 ( .ip1(\x[117][12] ), .ip2(n24450), .op(n22741) );
  nand2_1 U26713 ( .ip1(n22748), .ip2(n22741), .op(n22593) );
  nand2_1 U26714 ( .ip1(n24332), .ip2(\x[117][13] ), .op(n22742) );
  inv_1 U26715 ( .ip(n22742), .op(n22592) );
  inv_1 U26716 ( .ip(n22589), .op(n22591) );
  nand2_1 U26717 ( .ip1(\x[117][14] ), .ip2(n24230), .op(n22590) );
  nand2_1 U26718 ( .ip1(n22591), .ip2(n22590), .op(n22751) );
  not_ab_or_c_or_d U26719 ( .ip1(n22745), .ip2(n22593), .ip3(n22592), .ip4(
        n22751), .op(n22594) );
  nor4_1 U26720 ( .ip1(n22597), .ip2(n22596), .ip3(n22595), .ip4(n22594), .op(
        n24620) );
  inv_1 U26721 ( .ip(\x[120][12] ), .op(n22632) );
  and2_1 U26722 ( .ip1(n23146), .ip2(\x[120][10] ), .op(n22624) );
  inv_1 U26723 ( .ip(\x[120][9] ), .op(n22622) );
  and2_1 U26724 ( .ip1(n23804), .ip2(\x[120][8] ), .op(n22619) );
  inv_1 U26725 ( .ip(\x[120][7] ), .op(n22617) );
  nor2_1 U26726 ( .ip1(sig_in[7]), .ip2(n22617), .op(n22614) );
  inv_1 U26727 ( .ip(\x[120][3] ), .op(n22604) );
  nor2_1 U26728 ( .ip1(\x[120][2] ), .ip2(n23659), .op(n22603) );
  inv_1 U26729 ( .ip(\x[120][1] ), .op(n22599) );
  nor2_1 U26730 ( .ip1(sig_in[1]), .ip2(n22599), .op(n22601) );
  inv_1 U26731 ( .ip(\x[120][0] ), .op(n22598) );
  not_ab_or_c_or_d U26732 ( .ip1(n24467), .ip2(n22599), .ip3(n23195), .ip4(
        n22598), .op(n22600) );
  not_ab_or_c_or_d U26733 ( .ip1(\x[120][2] ), .ip2(n24470), .ip3(n22601), 
        .ip4(n22600), .op(n22602) );
  not_ab_or_c_or_d U26734 ( .ip1(sig_in[3]), .ip2(n22604), .ip3(n22603), .ip4(
        n22602), .op(n22608) );
  nand2_1 U26735 ( .ip1(\x[120][5] ), .ip2(n24119), .op(n22606) );
  nand2_1 U26736 ( .ip1(\x[120][4] ), .ip2(n23721), .op(n22605) );
  nand2_1 U26737 ( .ip1(n22606), .ip2(n22605), .op(n22607) );
  not_ab_or_c_or_d U26738 ( .ip1(\x[120][3] ), .ip2(n24342), .ip3(n22608), 
        .ip4(n22607), .op(n22612) );
  nor2_1 U26739 ( .ip1(\x[120][6] ), .ip2(n23770), .op(n22611) );
  nor2_1 U26740 ( .ip1(\x[120][5] ), .ip2(n24350), .op(n22610) );
  not_ab_or_c_or_d U26741 ( .ip1(\x[120][5] ), .ip2(n24482), .ip3(\x[120][4] ), 
        .ip4(n24256), .op(n22609) );
  nor4_1 U26742 ( .ip1(n22612), .ip2(n22611), .ip3(n22610), .ip4(n22609), .op(
        n22613) );
  not_ab_or_c_or_d U26743 ( .ip1(\x[120][6] ), .ip2(n24485), .ip3(n22614), 
        .ip4(n22613), .op(n22616) );
  nor2_1 U26744 ( .ip1(\x[120][8] ), .ip2(n23971), .op(n22615) );
  not_ab_or_c_or_d U26745 ( .ip1(sig_in[7]), .ip2(n22617), .ip3(n22616), .ip4(
        n22615), .op(n22618) );
  not_ab_or_c_or_d U26746 ( .ip1(\x[120][9] ), .ip2(n23981), .ip3(n22619), 
        .ip4(n22618), .op(n22621) );
  nor2_1 U26747 ( .ip1(\x[120][10] ), .ip2(n23980), .op(n22620) );
  not_ab_or_c_or_d U26748 ( .ip1(sig_in[9]), .ip2(n22622), .ip3(n22621), .ip4(
        n22620), .op(n22623) );
  not_ab_or_c_or_d U26749 ( .ip1(\x[120][11] ), .ip2(n24456), .ip3(n22624), 
        .ip4(n22623), .op(n22626) );
  nor2_1 U26750 ( .ip1(\x[120][11] ), .ip2(n24456), .op(n22625) );
  nor2_1 U26751 ( .ip1(n22626), .ip2(n22625), .op(n22627) );
  or2_1 U26752 ( .ip1(\x[120][12] ), .ip2(n22627), .op(n22629) );
  or2_1 U26753 ( .ip1(n24449), .ip2(n22627), .op(n22628) );
  nand2_1 U26754 ( .ip1(n22629), .ip2(n22628), .op(n22631) );
  nor2_1 U26755 ( .ip1(\x[120][13] ), .ip2(n24081), .op(n22630) );
  not_ab_or_c_or_d U26756 ( .ip1(sig_in[12]), .ip2(n22632), .ip3(n22631), 
        .ip4(n22630), .op(n22633) );
  nor2_1 U26757 ( .ip1(\x[120][15] ), .ip2(n24090), .op(n22634) );
  not_ab_or_c_or_d U26758 ( .ip1(\x[120][14] ), .ip2(n24230), .ip3(n22633), 
        .ip4(n22634), .op(n22680) );
  nand2_1 U26759 ( .ip1(\x[120][13] ), .ip2(n24235), .op(n22679) );
  nor3_1 U26760 ( .ip1(n22634), .ip2(\x[120][14] ), .ip3(n24382), .op(n22678)
         );
  nor2_1 U26761 ( .ip1(\x[119][15] ), .ip2(n24090), .op(n22733) );
  nor2_1 U26762 ( .ip1(\x[119][13] ), .ip2(n24081), .op(n22635) );
  or2_1 U26763 ( .ip1(sig_in[12]), .ip2(n22635), .op(n22638) );
  inv_1 U26764 ( .ip(\x[119][12] ), .op(n22636) );
  or2_1 U26765 ( .ip1(n22636), .ip2(n22635), .op(n22637) );
  nand2_1 U26766 ( .ip1(n22638), .ip2(n22637), .op(n22728) );
  and2_1 U26767 ( .ip1(n23146), .ip2(\x[119][10] ), .op(n22667) );
  inv_1 U26768 ( .ip(\x[119][9] ), .op(n22665) );
  and2_1 U26769 ( .ip1(n23804), .ip2(\x[119][8] ), .op(n22662) );
  inv_1 U26770 ( .ip(\x[119][7] ), .op(n22660) );
  nor2_1 U26771 ( .ip1(sig_in[7]), .ip2(n22660), .op(n22657) );
  inv_1 U26772 ( .ip(\x[119][5] ), .op(n22655) );
  nor2_1 U26773 ( .ip1(sig_in[5]), .ip2(n22655), .op(n22652) );
  inv_1 U26774 ( .ip(\x[119][3] ), .op(n22650) );
  and2_1 U26775 ( .ip1(n24335), .ip2(\x[119][2] ), .op(n22647) );
  inv_1 U26776 ( .ip(\x[119][1] ), .op(n22640) );
  inv_1 U26777 ( .ip(\x[119][0] ), .op(n22639) );
  not_ab_or_c_or_d U26778 ( .ip1(n24464), .ip2(n22640), .ip3(n23195), .ip4(
        n22639), .op(n22641) );
  or2_1 U26779 ( .ip1(\x[119][1] ), .ip2(n22641), .op(n22643) );
  or2_1 U26780 ( .ip1(n20652), .ip2(n22641), .op(n22642) );
  nand2_1 U26781 ( .ip1(n22643), .ip2(n22642), .op(n22645) );
  nor2_1 U26782 ( .ip1(\x[119][2] ), .ip2(n23659), .op(n22644) );
  nor2_1 U26783 ( .ip1(n22645), .ip2(n22644), .op(n22646) );
  not_ab_or_c_or_d U26784 ( .ip1(\x[119][3] ), .ip2(n24342), .ip3(n22647), 
        .ip4(n22646), .op(n22649) );
  nor2_1 U26785 ( .ip1(\x[119][4] ), .ip2(n24256), .op(n22648) );
  not_ab_or_c_or_d U26786 ( .ip1(sig_in[3]), .ip2(n22650), .ip3(n22649), .ip4(
        n22648), .op(n22651) );
  not_ab_or_c_or_d U26787 ( .ip1(\x[119][4] ), .ip2(n23860), .ip3(n22652), 
        .ip4(n22651), .op(n22654) );
  nor2_1 U26788 ( .ip1(\x[119][6] ), .ip2(n23509), .op(n22653) );
  not_ab_or_c_or_d U26789 ( .ip1(sig_in[5]), .ip2(n22655), .ip3(n22654), .ip4(
        n22653), .op(n22656) );
  not_ab_or_c_or_d U26790 ( .ip1(\x[119][6] ), .ip2(n23770), .ip3(n22657), 
        .ip4(n22656), .op(n22659) );
  nor2_1 U26791 ( .ip1(\x[119][8] ), .ip2(n23971), .op(n22658) );
  not_ab_or_c_or_d U26792 ( .ip1(sig_in[7]), .ip2(n22660), .ip3(n22659), .ip4(
        n22658), .op(n22661) );
  not_ab_or_c_or_d U26793 ( .ip1(\x[119][9] ), .ip2(n24043), .ip3(n22662), 
        .ip4(n22661), .op(n22664) );
  nor2_1 U26794 ( .ip1(\x[119][10] ), .ip2(n24370), .op(n22663) );
  not_ab_or_c_or_d U26795 ( .ip1(sig_in[9]), .ip2(n22665), .ip3(n22664), .ip4(
        n22663), .op(n22666) );
  not_ab_or_c_or_d U26796 ( .ip1(\x[119][11] ), .ip2(n24456), .ip3(n22667), 
        .ip4(n22666), .op(n22669) );
  nor2_1 U26797 ( .ip1(\x[119][11] ), .ip2(n21793), .op(n22668) );
  nor2_1 U26798 ( .ip1(n22669), .ip2(n22668), .op(n22726) );
  inv_1 U26799 ( .ip(\x[119][14] ), .op(n22672) );
  nor2_1 U26800 ( .ip1(sig_in[14]), .ip2(n22672), .op(n22730) );
  nand2_1 U26801 ( .ip1(\x[119][13] ), .ip2(n24235), .op(n22671) );
  nand2_1 U26802 ( .ip1(\x[119][12] ), .ip2(n24079), .op(n22670) );
  nand2_1 U26803 ( .ip1(n22671), .ip2(n22670), .op(n22727) );
  not_ab_or_c_or_d U26804 ( .ip1(n22728), .ip2(n22726), .ip3(n22730), .ip4(
        n22727), .op(n22675) );
  nand2_1 U26805 ( .ip1(sig_in[14]), .ip2(n22672), .op(n22674) );
  nand2_1 U26806 ( .ip1(\x[119][15] ), .ip2(n24180), .op(n22673) );
  nand2_1 U26807 ( .ip1(n22674), .ip2(n22673), .op(n22735) );
  nor2_1 U26808 ( .ip1(n22675), .ip2(n22735), .op(n22676) );
  ab_or_c_or_d U26809 ( .ip1(\x[120][15] ), .ip2(n24180), .ip3(n22733), .ip4(
        n22676), .op(n22677) );
  not_ab_or_c_or_d U26810 ( .ip1(n22680), .ip2(n22679), .ip3(n22678), .ip4(
        n22677), .op(n27300) );
  and2_1 U26811 ( .ip1(n24332), .ip2(\x[118][13] ), .op(n22681) );
  nor2_1 U26812 ( .ip1(\x[118][15] ), .ip2(n24090), .op(n22686) );
  not_ab_or_c_or_d U26813 ( .ip1(\x[118][14] ), .ip2(n24230), .ip3(n22681), 
        .ip4(n22686), .op(n22757) );
  nand2_1 U26814 ( .ip1(\x[118][12] ), .ip2(n24450), .op(n22682) );
  nand2_1 U26815 ( .ip1(n22757), .ip2(n22682), .op(n22753) );
  nor2_1 U26816 ( .ip1(\x[118][14] ), .ip2(n24382), .op(n22683) );
  or2_1 U26817 ( .ip1(\x[118][15] ), .ip2(n22683), .op(n22685) );
  or2_1 U26818 ( .ip1(n24329), .ip2(n22683), .op(n22684) );
  nand2_1 U26819 ( .ip1(n22685), .ip2(n22684), .op(n22724) );
  or2_1 U26820 ( .ip1(n22686), .ip2(n22724), .op(n22758) );
  nor2_1 U26821 ( .ip1(\x[118][9] ), .ip2(n24269), .op(n22711) );
  inv_1 U26822 ( .ip(\x[118][8] ), .op(n22687) );
  nor3_1 U26823 ( .ip1(sig_in[8]), .ip2(n22711), .ip3(n22687), .op(n22714) );
  and2_1 U26824 ( .ip1(n24461), .ip2(\x[118][7] ), .op(n22708) );
  inv_1 U26825 ( .ip(\x[118][5] ), .op(n22706) );
  inv_1 U26826 ( .ip(\x[118][4] ), .op(n22698) );
  nor2_1 U26827 ( .ip1(n24462), .ip2(n22698), .op(n22696) );
  inv_1 U26828 ( .ip(\x[118][3] ), .op(n22694) );
  inv_1 U26829 ( .ip(\x[118][1] ), .op(n22689) );
  nor2_1 U26830 ( .ip1(sig_in[1]), .ip2(n22689), .op(n22691) );
  inv_1 U26831 ( .ip(\x[118][0] ), .op(n22688) );
  not_ab_or_c_or_d U26832 ( .ip1(n24467), .ip2(n22689), .ip3(n23195), .ip4(
        n22688), .op(n22690) );
  not_ab_or_c_or_d U26833 ( .ip1(\x[118][2] ), .ip2(n24470), .ip3(n22691), 
        .ip4(n22690), .op(n22693) );
  nor2_1 U26834 ( .ip1(\x[118][2] ), .ip2(n23717), .op(n22692) );
  not_ab_or_c_or_d U26835 ( .ip1(sig_in[3]), .ip2(n22694), .ip3(n22693), .ip4(
        n22692), .op(n22695) );
  not_ab_or_c_or_d U26836 ( .ip1(\x[118][3] ), .ip2(n24342), .ip3(n22696), 
        .ip4(n22695), .op(n22697) );
  or2_1 U26837 ( .ip1(sig_in[4]), .ip2(n22697), .op(n22700) );
  or2_1 U26838 ( .ip1(n22698), .ip2(n22697), .op(n22699) );
  nand2_1 U26839 ( .ip1(n22700), .ip2(n22699), .op(n22701) );
  or2_1 U26840 ( .ip1(\x[118][5] ), .ip2(n22701), .op(n22703) );
  or2_1 U26841 ( .ip1(n23600), .ip2(n22701), .op(n22702) );
  nand2_1 U26842 ( .ip1(n22703), .ip2(n22702), .op(n22705) );
  nor2_1 U26843 ( .ip1(\x[118][6] ), .ip2(n24355), .op(n22704) );
  not_ab_or_c_or_d U26844 ( .ip1(n22833), .ip2(n22706), .ip3(n22705), .ip4(
        n22704), .op(n22707) );
  not_ab_or_c_or_d U26845 ( .ip1(\x[118][6] ), .ip2(n23509), .ip3(n22708), 
        .ip4(n22707), .op(n22712) );
  nor2_1 U26846 ( .ip1(\x[118][7] ), .ip2(n24492), .op(n22710) );
  nor2_1 U26847 ( .ip1(\x[118][8] ), .ip2(n24100), .op(n22709) );
  nor4_1 U26848 ( .ip1(n22712), .ip2(n22711), .ip3(n22710), .ip4(n22709), .op(
        n22713) );
  not_ab_or_c_or_d U26849 ( .ip1(\x[118][10] ), .ip2(n23980), .ip3(n22714), 
        .ip4(n22713), .op(n22718) );
  nand2_1 U26850 ( .ip1(\x[118][9] ), .ip2(n24043), .op(n22717) );
  nor2_1 U26851 ( .ip1(\x[118][10] ), .ip2(n23980), .op(n22716) );
  nor2_1 U26852 ( .ip1(\x[118][11] ), .ip2(n21793), .op(n22715) );
  not_ab_or_c_or_d U26853 ( .ip1(n22718), .ip2(n22717), .ip3(n22716), .ip4(
        n22715), .op(n22719) );
  or2_1 U26854 ( .ip1(\x[118][11] ), .ip2(n22719), .op(n22721) );
  or2_1 U26855 ( .ip1(n24136), .ip2(n22719), .op(n22720) );
  nand2_1 U26856 ( .ip1(n22721), .ip2(n22720), .op(n22754) );
  nor2_1 U26857 ( .ip1(\x[118][13] ), .ip2(n24081), .op(n22723) );
  nor2_1 U26858 ( .ip1(\x[118][12] ), .ip2(n24079), .op(n22722) );
  or2_1 U26859 ( .ip1(n22723), .ip2(n22722), .op(n22756) );
  inv_1 U26860 ( .ip(n22724), .op(n22725) );
  nor3_1 U26861 ( .ip1(n22754), .ip2(n22756), .ip3(n22725), .op(n22739) );
  or2_1 U26862 ( .ip1(n22727), .ip2(n22726), .op(n22729) );
  nand2_1 U26863 ( .ip1(n22729), .ip2(n22728), .op(n22732) );
  nor2_1 U26864 ( .ip1(n22730), .ip2(n22733), .op(n22731) );
  nand2_1 U26865 ( .ip1(n22732), .ip2(n22731), .op(n22737) );
  inv_1 U26866 ( .ip(n22733), .op(n22734) );
  nand2_1 U26867 ( .ip1(n22735), .ip2(n22734), .op(n22736) );
  nand2_1 U26868 ( .ip1(n22737), .ip2(n22736), .op(n22738) );
  not_ab_or_c_or_d U26869 ( .ip1(n22753), .ip2(n22758), .ip3(n22739), .ip4(
        n22738), .op(n27299) );
  nor2_1 U26870 ( .ip1(n27300), .ip2(n27299), .op(n24626) );
  inv_1 U26871 ( .ip(n22740), .op(n22747) );
  or2_1 U26872 ( .ip1(n22741), .ip2(n22747), .op(n22744) );
  or2_1 U26873 ( .ip1(n22742), .ip2(n22747), .op(n22743) );
  nand2_1 U26874 ( .ip1(n22744), .ip2(n22743), .op(n22750) );
  inv_1 U26875 ( .ip(n22745), .op(n22746) );
  nor3_1 U26876 ( .ip1(n22748), .ip2(n22747), .ip3(n22746), .op(n22749) );
  not_ab_or_c_or_d U26877 ( .ip1(n22752), .ip2(n22751), .ip3(n22750), .ip4(
        n22749), .op(n22761) );
  inv_1 U26878 ( .ip(n22753), .op(n22755) );
  nand2_1 U26879 ( .ip1(n22755), .ip2(n22754), .op(n22760) );
  nand2_1 U26880 ( .ip1(n22757), .ip2(n22756), .op(n22759) );
  nand4_1 U26881 ( .ip1(n22761), .ip2(n22760), .ip3(n22759), .ip4(n22758), 
        .op(n24628) );
  nand2_1 U26882 ( .ip1(n24626), .ip2(n24628), .op(n24621) );
  nor2_1 U26883 ( .ip1(n24620), .ip2(n24621), .op(n24623) );
  inv_1 U26884 ( .ip(n22762), .op(n22763) );
  nor2_1 U26885 ( .ip1(n22764), .ip2(n22763), .op(n22771) );
  inv_1 U26886 ( .ip(n22765), .op(n22767) );
  nor2_1 U26887 ( .ip1(n22767), .ip2(n22766), .op(n22768) );
  nor2_1 U26888 ( .ip1(n22769), .ip2(n22768), .op(n22770) );
  not_ab_or_c_or_d U26889 ( .ip1(n22773), .ip2(n22772), .ip3(n22771), .ip4(
        n22770), .op(n22777) );
  inv_1 U26890 ( .ip(n22774), .op(n22776) );
  nand3_1 U26891 ( .ip1(n22777), .ip2(n22776), .ip3(n22775), .op(n24625) );
  nand2_1 U26892 ( .ip1(n24623), .ip2(n24625), .op(n24640) );
  nor2_1 U26893 ( .ip1(n24639), .ip2(n24640), .op(n24636) );
  or2_1 U26894 ( .ip1(n22779), .ip2(n22778), .op(n22793) );
  inv_1 U26895 ( .ip(n22780), .op(n22787) );
  inv_1 U26896 ( .ip(n22781), .op(n22783) );
  nor3_1 U26897 ( .ip1(n22784), .ip2(n22783), .ip3(n22782), .op(n22786) );
  not_ab_or_c_or_d U26898 ( .ip1(n22788), .ip2(n22787), .ip3(n22786), .ip4(
        n22785), .op(n22792) );
  or2_1 U26899 ( .ip1(n22790), .ip2(n22789), .op(n22791) );
  nand3_1 U26900 ( .ip1(n22793), .ip2(n22792), .ip3(n22791), .op(n24638) );
  nand2_1 U26901 ( .ip1(n24636), .ip2(n24638), .op(n27371) );
  nor4_1 U26902 ( .ip1(n24569), .ip2(n24571), .ip3(n27142), .ip4(n27371), .op(
        n27288) );
  nor2_1 U26903 ( .ip1(\x[2][9] ), .ip2(n24164), .op(n22818) );
  inv_1 U26904 ( .ip(\x[2][8] ), .op(n22794) );
  nor3_1 U26905 ( .ip1(sig_in[8]), .ip2(n22818), .ip3(n22794), .op(n22822) );
  nor2_1 U26906 ( .ip1(\x[2][7] ), .ip2(n24044), .op(n22820) );
  nor2_1 U26907 ( .ip1(\x[2][8] ), .ip2(n23971), .op(n22819) );
  and2_1 U26908 ( .ip1(n23770), .ip2(\x[2][6] ), .op(n22811) );
  inv_1 U26909 ( .ip(\x[2][3] ), .op(n22804) );
  and2_1 U26910 ( .ip1(n24107), .ip2(\x[2][2] ), .op(n22801) );
  nand2_1 U26911 ( .ip1(\x[2][1] ), .ip2(n21685), .op(n22799) );
  nand2_1 U26912 ( .ip1(\x[2][0] ), .ip2(n24143), .op(n22798) );
  nor2_1 U26913 ( .ip1(\x[2][2] ), .ip2(n23659), .op(n22797) );
  nor2_1 U26914 ( .ip1(\x[2][1] ), .ip2(n20652), .op(n22796) );
  not_ab_or_c_or_d U26915 ( .ip1(n22799), .ip2(n22798), .ip3(n22797), .ip4(
        n22796), .op(n22800) );
  not_ab_or_c_or_d U26916 ( .ip1(\x[2][3] ), .ip2(n24342), .ip3(n22801), .ip4(
        n22800), .op(n22803) );
  nor2_1 U26917 ( .ip1(\x[2][4] ), .ip2(n23860), .op(n22802) );
  not_ab_or_c_or_d U26918 ( .ip1(n24251), .ip2(n22804), .ip3(n22803), .ip4(
        n22802), .op(n22805) );
  or2_1 U26919 ( .ip1(\x[2][4] ), .ip2(n22805), .op(n22807) );
  or2_1 U26920 ( .ip1(n23860), .ip2(n22805), .op(n22806) );
  nand2_1 U26921 ( .ip1(n22807), .ip2(n22806), .op(n22809) );
  nor2_1 U26922 ( .ip1(\x[2][5] ), .ip2(n24350), .op(n22808) );
  nor2_1 U26923 ( .ip1(n22809), .ip2(n22808), .op(n22810) );
  not_ab_or_c_or_d U26924 ( .ip1(\x[2][5] ), .ip2(n23600), .ip3(n22811), .ip4(
        n22810), .op(n22813) );
  nor2_1 U26925 ( .ip1(\x[2][6] ), .ip2(n24355), .op(n22812) );
  nor2_1 U26926 ( .ip1(n22813), .ip2(n22812), .op(n22814) );
  or2_1 U26927 ( .ip1(\x[2][7] ), .ip2(n22814), .op(n22816) );
  or2_1 U26928 ( .ip1(n24142), .ip2(n22814), .op(n22815) );
  nand2_1 U26929 ( .ip1(n22816), .ip2(n22815), .op(n22817) );
  nor4_1 U26930 ( .ip1(n22820), .ip2(n22819), .ip3(n22818), .ip4(n22817), .op(
        n22821) );
  not_ab_or_c_or_d U26931 ( .ip1(\x[2][9] ), .ip2(n24455), .ip3(n22822), .ip4(
        n22821), .op(n22826) );
  nand2_1 U26932 ( .ip1(\x[2][10] ), .ip2(n23146), .op(n22825) );
  nor2_1 U26933 ( .ip1(\x[2][10] ), .ip2(n23980), .op(n22824) );
  nor2_1 U26934 ( .ip1(\x[2][11] ), .ip2(n21793), .op(n22823) );
  not_ab_or_c_or_d U26935 ( .ip1(n22826), .ip2(n22825), .ip3(n22824), .ip4(
        n22823), .op(n22827) );
  or2_1 U26936 ( .ip1(\x[2][11] ), .ip2(n22827), .op(n22829) );
  or2_1 U26937 ( .ip1(n24136), .ip2(n22827), .op(n22828) );
  nand2_1 U26938 ( .ip1(n22829), .ip2(n22828), .op(n23626) );
  and2_1 U26939 ( .ip1(n23895), .ip2(\x[2][13] ), .op(n22832) );
  inv_1 U26940 ( .ip(\x[2][15] ), .op(n22878) );
  nand2_1 U26941 ( .ip1(sig_in[15]), .ip2(n22878), .op(n22831) );
  nand2_1 U26942 ( .ip1(\x[2][14] ), .ip2(n24327), .op(n22830) );
  nand2_1 U26943 ( .ip1(n22831), .ip2(n22830), .op(n22877) );
  not_ab_or_c_or_d U26944 ( .ip1(\x[2][12] ), .ip2(n24449), .ip3(n22832), 
        .ip4(n22877), .op(n23624) );
  inv_1 U26945 ( .ip(\x[1][12] ), .op(n22872) );
  nor2_1 U26946 ( .ip1(\x[1][11] ), .ip2(n24456), .op(n22863) );
  nor2_1 U26947 ( .ip1(\x[1][9] ), .ip2(n24043), .op(n22862) );
  nor2_1 U26948 ( .ip1(\x[1][10] ), .ip2(n24370), .op(n22861) );
  and2_1 U26949 ( .ip1(n23804), .ip2(\x[1][8] ), .op(n22855) );
  inv_1 U26950 ( .ip(\x[1][6] ), .op(n22853) );
  inv_1 U26951 ( .ip(\x[1][5] ), .op(n22845) );
  nor2_1 U26952 ( .ip1(n22845), .ip2(n22833), .op(n22847) );
  nor2_1 U26953 ( .ip1(\x[1][4] ), .ip2(n24347), .op(n22844) );
  and2_1 U26954 ( .ip1(n23721), .ip2(\x[1][4] ), .op(n22842) );
  inv_1 U26955 ( .ip(\x[1][3] ), .op(n22840) );
  inv_1 U26956 ( .ip(\x[1][1] ), .op(n22835) );
  nor2_1 U26957 ( .ip1(sig_in[1]), .ip2(n22835), .op(n22837) );
  inv_1 U26958 ( .ip(\x[1][0] ), .op(n22834) );
  not_ab_or_c_or_d U26959 ( .ip1(n24464), .ip2(n22835), .ip3(n23195), .ip4(
        n22834), .op(n22836) );
  not_ab_or_c_or_d U26960 ( .ip1(\x[1][2] ), .ip2(n24470), .ip3(n22837), .ip4(
        n22836), .op(n22839) );
  nor2_1 U26961 ( .ip1(\x[1][2] ), .ip2(n24107), .op(n22838) );
  not_ab_or_c_or_d U26962 ( .ip1(n23251), .ip2(n22840), .ip3(n22839), .ip4(
        n22838), .op(n22841) );
  not_ab_or_c_or_d U26963 ( .ip1(\x[1][3] ), .ip2(n22795), .ip3(n22842), .ip4(
        n22841), .op(n22843) );
  not_ab_or_c_or_d U26964 ( .ip1(n22833), .ip2(n22845), .ip3(n22844), .ip4(
        n22843), .op(n22846) );
  or2_1 U26965 ( .ip1(n22847), .ip2(n22846), .op(n22848) );
  or2_1 U26966 ( .ip1(\x[1][6] ), .ip2(n22848), .op(n22850) );
  or2_1 U26967 ( .ip1(n23509), .ip2(n22848), .op(n22849) );
  nand2_1 U26968 ( .ip1(n22850), .ip2(n22849), .op(n22852) );
  nor2_1 U26969 ( .ip1(\x[1][7] ), .ip2(n24492), .op(n22851) );
  not_ab_or_c_or_d U26970 ( .ip1(sig_in[6]), .ip2(n22853), .ip3(n22852), .ip4(
        n22851), .op(n22854) );
  not_ab_or_c_or_d U26971 ( .ip1(\x[1][7] ), .ip2(n24142), .ip3(n22855), .ip4(
        n22854), .op(n22857) );
  nor2_1 U26972 ( .ip1(n24358), .ip2(\x[1][8] ), .op(n22856) );
  nor2_1 U26973 ( .ip1(n22857), .ip2(n22856), .op(n22859) );
  and2_1 U26974 ( .ip1(n23981), .ip2(\x[1][9] ), .op(n22858) );
  nor2_1 U26975 ( .ip1(n22859), .ip2(n22858), .op(n22860) );
  nor4_1 U26976 ( .ip1(n22863), .ip2(n22862), .ip3(n22861), .ip4(n22860), .op(
        n22869) );
  nand2_1 U26977 ( .ip1(n24456), .ip2(\x[1][11] ), .op(n22867) );
  inv_1 U26978 ( .ip(n22863), .op(n22864) );
  nand3_1 U26979 ( .ip1(\x[1][10] ), .ip2(n23980), .ip3(n22864), .op(n22866)
         );
  nand2_1 U26980 ( .ip1(\x[1][13] ), .ip2(n24081), .op(n22865) );
  nand3_1 U26981 ( .ip1(n22867), .ip2(n22866), .ip3(n22865), .op(n22868) );
  not_ab_or_c_or_d U26982 ( .ip1(\x[1][12] ), .ip2(n24449), .ip3(n22869), 
        .ip4(n22868), .op(n22871) );
  nor2_1 U26983 ( .ip1(\x[1][13] ), .ip2(n24376), .op(n22870) );
  not_ab_or_c_or_d U26984 ( .ip1(sig_in[12]), .ip2(n22872), .ip3(n22871), 
        .ip4(n22870), .op(n22874) );
  nor2_1 U26985 ( .ip1(\x[1][15] ), .ip2(n24090), .op(n22873) );
  nor3_1 U26986 ( .ip1(\x[1][14] ), .ip2(n22874), .ip3(n22873), .op(n22876) );
  not_ab_or_c_or_d U26987 ( .ip1(n22874), .ip2(\x[1][14] ), .ip3(n22873), 
        .ip4(n23938), .op(n22875) );
  nor2_1 U26988 ( .ip1(n22876), .ip2(n22875), .op(n24515) );
  nand2_1 U26989 ( .ip1(n23143), .ip2(\x[1][15] ), .op(n24514) );
  and2_1 U26990 ( .ip1(n24515), .ip2(n24514), .op(n22886) );
  inv_1 U26991 ( .ip(n22877), .op(n22879) );
  nor2_1 U26992 ( .ip1(sig_in[15]), .ip2(n22878), .op(n22880) );
  nor2_1 U26993 ( .ip1(n22879), .ip2(n22880), .op(n23621) );
  or2_1 U26994 ( .ip1(n24233), .ip2(\x[2][12] ), .op(n22883) );
  inv_1 U26995 ( .ip(\x[2][14] ), .op(n22882) );
  nor2_1 U26996 ( .ip1(\x[2][13] ), .ip2(n24376), .op(n22881) );
  not_ab_or_c_or_d U26997 ( .ip1(sig_in[14]), .ip2(n22882), .ip3(n22881), 
        .ip4(n22880), .op(n23622) );
  nand2_1 U26998 ( .ip1(n22883), .ip2(n23622), .op(n23625) );
  inv_1 U26999 ( .ip(n23625), .op(n22884) );
  nor2_1 U27000 ( .ip1(n23621), .ip2(n22884), .op(n22885) );
  not_ab_or_c_or_d U27001 ( .ip1(n23626), .ip2(n23624), .ip3(n22886), .ip4(
        n22885), .op(n24758) );
  inv_1 U27002 ( .ip(\x[4][11] ), .op(n22919) );
  nor2_1 U27003 ( .ip1(n22919), .ip2(n17981), .op(n22921) );
  nor2_1 U27004 ( .ip1(\x[4][10] ), .ip2(n23980), .op(n22918) );
  and2_1 U27005 ( .ip1(n24451), .ip2(\x[4][10] ), .op(n22916) );
  inv_1 U27006 ( .ip(\x[4][9] ), .op(n22914) );
  nor2_1 U27007 ( .ip1(\x[4][8] ), .ip2(n24100), .op(n22913) );
  inv_1 U27008 ( .ip(\x[4][7] ), .op(n22908) );
  and2_1 U27009 ( .ip1(n24335), .ip2(\x[4][2] ), .op(n22895) );
  inv_1 U27010 ( .ip(\x[4][1] ), .op(n22888) );
  inv_1 U27011 ( .ip(\x[4][0] ), .op(n22887) );
  not_ab_or_c_or_d U27012 ( .ip1(n24467), .ip2(n22888), .ip3(n23195), .ip4(
        n22887), .op(n22889) );
  or2_1 U27013 ( .ip1(\x[4][1] ), .ip2(n22889), .op(n22891) );
  or2_1 U27014 ( .ip1(n20652), .ip2(n22889), .op(n22890) );
  nand2_1 U27015 ( .ip1(n22891), .ip2(n22890), .op(n22893) );
  nor2_1 U27016 ( .ip1(\x[4][2] ), .ip2(n23659), .op(n22892) );
  nor2_1 U27017 ( .ip1(n22893), .ip2(n22892), .op(n22894) );
  not_ab_or_c_or_d U27018 ( .ip1(\x[4][3] ), .ip2(n24476), .ip3(n22895), .ip4(
        n22894), .op(n22898) );
  nor2_1 U27019 ( .ip1(\x[4][5] ), .ip2(n24350), .op(n22899) );
  nor2_1 U27020 ( .ip1(\x[4][4] ), .ip2(n23721), .op(n22897) );
  nor2_1 U27021 ( .ip1(\x[4][3] ), .ip2(n24342), .op(n22896) );
  nor4_1 U27022 ( .ip1(n22898), .ip2(n22899), .ip3(n22897), .ip4(n22896), .op(
        n22905) );
  nand2_1 U27023 ( .ip1(n23600), .ip2(\x[4][5] ), .op(n22903) );
  inv_1 U27024 ( .ip(n22899), .op(n22900) );
  nand3_1 U27025 ( .ip1(\x[4][4] ), .ip2(n23721), .ip3(n22900), .op(n22902) );
  nand2_1 U27026 ( .ip1(\x[4][7] ), .ip2(n24044), .op(n22901) );
  nand3_1 U27027 ( .ip1(n22903), .ip2(n22902), .ip3(n22901), .op(n22904) );
  not_ab_or_c_or_d U27028 ( .ip1(\x[4][6] ), .ip2(n23770), .ip3(n22905), .ip4(
        n22904), .op(n22907) );
  not_ab_or_c_or_d U27029 ( .ip1(\x[4][7] ), .ip2(n24461), .ip3(\x[4][6] ), 
        .ip4(n23770), .op(n22906) );
  not_ab_or_c_or_d U27030 ( .ip1(sig_in[7]), .ip2(n22908), .ip3(n22907), .ip4(
        n22906), .op(n22909) );
  or2_1 U27031 ( .ip1(\x[4][8] ), .ip2(n22909), .op(n22911) );
  or2_1 U27032 ( .ip1(n24100), .ip2(n22909), .op(n22910) );
  nand2_1 U27033 ( .ip1(n22911), .ip2(n22910), .op(n22912) );
  not_ab_or_c_or_d U27034 ( .ip1(sig_in[9]), .ip2(n22914), .ip3(n22913), .ip4(
        n22912), .op(n22915) );
  not_ab_or_c_or_d U27035 ( .ip1(\x[4][9] ), .ip2(n24455), .ip3(n22916), .ip4(
        n22915), .op(n22917) );
  not_ab_or_c_or_d U27036 ( .ip1(sig_in[11]), .ip2(n22919), .ip3(n22918), 
        .ip4(n22917), .op(n22920) );
  or2_1 U27037 ( .ip1(n22921), .ip2(n22920), .op(n23638) );
  and2_1 U27038 ( .ip1(n24186), .ip2(\x[4][15] ), .op(n22977) );
  nor2_1 U27039 ( .ip1(\x[4][14] ), .ip2(n23938), .op(n22924) );
  nor2_1 U27040 ( .ip1(\x[4][13] ), .ip2(n24137), .op(n22923) );
  nor2_1 U27041 ( .ip1(\x[4][12] ), .ip2(n24233), .op(n22922) );
  nor4_1 U27042 ( .ip1(n22977), .ip2(n22924), .ip3(n22923), .ip4(n22922), .op(
        n23640) );
  nor2_1 U27043 ( .ip1(\x[5][14] ), .ip2(n24185), .op(n22925) );
  or2_1 U27044 ( .ip1(\x[5][15] ), .ip2(n22925), .op(n22927) );
  or2_1 U27045 ( .ip1(n24384), .ip2(n22925), .op(n22926) );
  nand2_1 U27046 ( .ip1(n22927), .ip2(n22926), .op(n22994) );
  nor2_1 U27047 ( .ip1(\x[5][15] ), .ip2(n24329), .op(n23043) );
  or2_1 U27048 ( .ip1(n22994), .ip2(n23043), .op(n22973) );
  and2_1 U27049 ( .ip1(n23895), .ip2(\x[5][13] ), .op(n22928) );
  or2_1 U27050 ( .ip1(\x[5][14] ), .ip2(n22928), .op(n22930) );
  or2_1 U27051 ( .ip1(n24327), .ip2(n22928), .op(n22929) );
  nand2_1 U27052 ( .ip1(n22930), .ip2(n22929), .op(n22989) );
  nor2_1 U27053 ( .ip1(\x[5][13] ), .ip2(n24137), .op(n22931) );
  or2_1 U27054 ( .ip1(sig_in[12]), .ip2(n22931), .op(n22934) );
  inv_1 U27055 ( .ip(\x[5][12] ), .op(n22932) );
  or2_1 U27056 ( .ip1(n22932), .ip2(n22931), .op(n22933) );
  nand2_1 U27057 ( .ip1(n22934), .ip2(n22933), .op(n22993) );
  inv_1 U27058 ( .ip(\x[5][9] ), .op(n22959) );
  and2_1 U27059 ( .ip1(n24461), .ip2(\x[5][7] ), .op(n22951) );
  inv_1 U27060 ( .ip(n24342), .op(n23251) );
  inv_1 U27061 ( .ip(\x[5][3] ), .op(n22941) );
  nor2_1 U27062 ( .ip1(\x[5][2] ), .ip2(n23717), .op(n22940) );
  inv_1 U27063 ( .ip(\x[5][1] ), .op(n22936) );
  nor2_1 U27064 ( .ip1(sig_in[1]), .ip2(n22936), .op(n22938) );
  inv_1 U27065 ( .ip(\x[5][0] ), .op(n22935) );
  not_ab_or_c_or_d U27066 ( .ip1(n24467), .ip2(n22936), .ip3(n23195), .ip4(
        n22935), .op(n22937) );
  not_ab_or_c_or_d U27067 ( .ip1(\x[5][2] ), .ip2(n24470), .ip3(n22938), .ip4(
        n22937), .op(n22939) );
  not_ab_or_c_or_d U27068 ( .ip1(n23251), .ip2(n22941), .ip3(n22940), .ip4(
        n22939), .op(n22945) );
  nand2_1 U27069 ( .ip1(\x[5][5] ), .ip2(n24119), .op(n22943) );
  nand2_1 U27070 ( .ip1(\x[5][4] ), .ip2(n23721), .op(n22942) );
  nand2_1 U27071 ( .ip1(n22943), .ip2(n22942), .op(n22944) );
  not_ab_or_c_or_d U27072 ( .ip1(\x[5][3] ), .ip2(n24342), .ip3(n22945), .ip4(
        n22944), .op(n22949) );
  nor2_1 U27073 ( .ip1(\x[5][5] ), .ip2(n24350), .op(n22948) );
  nor2_1 U27074 ( .ip1(\x[5][6] ), .ip2(n24355), .op(n22947) );
  not_ab_or_c_or_d U27075 ( .ip1(\x[5][5] ), .ip2(n23600), .ip3(\x[5][4] ), 
        .ip4(n24256), .op(n22946) );
  nor4_1 U27076 ( .ip1(n22949), .ip2(n22948), .ip3(n22947), .ip4(n22946), .op(
        n22950) );
  not_ab_or_c_or_d U27077 ( .ip1(\x[5][6] ), .ip2(n24045), .ip3(n22951), .ip4(
        n22950), .op(n22953) );
  nor2_1 U27078 ( .ip1(\x[5][7] ), .ip2(n24492), .op(n22952) );
  nor2_1 U27079 ( .ip1(n22953), .ip2(n22952), .op(n22954) );
  or2_1 U27080 ( .ip1(\x[5][8] ), .ip2(n22954), .op(n22956) );
  or2_1 U27081 ( .ip1(n24100), .ip2(n22954), .op(n22955) );
  nand2_1 U27082 ( .ip1(n22956), .ip2(n22955), .op(n22958) );
  nor2_1 U27083 ( .ip1(\x[5][8] ), .ip2(n24100), .op(n22957) );
  not_ab_or_c_or_d U27084 ( .ip1(sig_in[9]), .ip2(n22959), .ip3(n22958), .ip4(
        n22957), .op(n22960) );
  or2_1 U27085 ( .ip1(\x[5][9] ), .ip2(n22960), .op(n22962) );
  or2_1 U27086 ( .ip1(n24164), .ip2(n22960), .op(n22961) );
  nand2_1 U27087 ( .ip1(n22962), .ip2(n22961), .op(n22983) );
  nand2_1 U27088 ( .ip1(\x[5][10] ), .ip2(n24370), .op(n22981) );
  nand2_1 U27089 ( .ip1(n22983), .ip2(n22981), .op(n22967) );
  nor2_1 U27090 ( .ip1(\x[5][11] ), .ip2(n21793), .op(n22986) );
  or2_1 U27091 ( .ip1(sig_in[10]), .ip2(n22986), .op(n22965) );
  inv_1 U27092 ( .ip(\x[5][10] ), .op(n22963) );
  or2_1 U27093 ( .ip1(n22963), .ip2(n22986), .op(n22964) );
  nand2_1 U27094 ( .ip1(n22965), .ip2(n22964), .op(n22966) );
  nand2_1 U27095 ( .ip1(n22967), .ip2(n22966), .op(n22968) );
  nand2_1 U27096 ( .ip1(\x[5][11] ), .ip2(n24239), .op(n22980) );
  nand2_1 U27097 ( .ip1(\x[5][12] ), .ip2(n24450), .op(n22988) );
  nand3_1 U27098 ( .ip1(n22968), .ip2(n22980), .ip3(n22988), .op(n22969) );
  nand2_1 U27099 ( .ip1(n22993), .ip2(n22969), .op(n22970) );
  nand2_1 U27100 ( .ip1(n22989), .ip2(n22970), .op(n22971) );
  or2_1 U27101 ( .ip1(n22971), .ip2(n23043), .op(n22972) );
  nand2_1 U27102 ( .ip1(n22973), .ip2(n22972), .op(n22979) );
  nor2_1 U27103 ( .ip1(\x[4][15] ), .ip2(n24090), .op(n23639) );
  nand2_1 U27104 ( .ip1(\x[4][13] ), .ip2(n24081), .op(n22975) );
  nand2_1 U27105 ( .ip1(\x[4][12] ), .ip2(n24233), .op(n22974) );
  nand2_1 U27106 ( .ip1(n22975), .ip2(n22974), .op(n22976) );
  not_ab_or_c_or_d U27107 ( .ip1(\x[4][14] ), .ip2(n23938), .ip3(n23639), 
        .ip4(n22976), .op(n23636) );
  nor2_1 U27108 ( .ip1(n22977), .ip2(n23636), .op(n22978) );
  not_ab_or_c_or_d U27109 ( .ip1(n23638), .ip2(n23640), .ip3(n22979), .ip4(
        n22978), .op(n24763) );
  nand2_1 U27110 ( .ip1(n22981), .ip2(n22980), .op(n22985) );
  nor2_1 U27111 ( .ip1(\x[5][10] ), .ip2(n23980), .op(n22982) );
  nor2_1 U27112 ( .ip1(n22983), .ip2(n22982), .op(n22984) );
  nor2_1 U27113 ( .ip1(n22985), .ip2(n22984), .op(n22987) );
  nor2_1 U27114 ( .ip1(n22987), .ip2(n22986), .op(n22992) );
  inv_1 U27115 ( .ip(n22988), .op(n22991) );
  inv_1 U27116 ( .ip(n22989), .op(n22990) );
  not_ab_or_c_or_d U27117 ( .ip1(n22993), .ip2(n22992), .ip3(n22991), .ip4(
        n22990), .op(n22996) );
  inv_1 U27118 ( .ip(n22994), .op(n22995) );
  nor2_1 U27119 ( .ip1(n22996), .ip2(n22995), .op(n23042) );
  nor2_1 U27120 ( .ip1(\x[6][15] ), .ip2(n24090), .op(n23001) );
  nand2_1 U27121 ( .ip1(n24384), .ip2(\x[6][15] ), .op(n23554) );
  inv_1 U27122 ( .ip(n23554), .op(n22997) );
  or2_1 U27123 ( .ip1(sig_in[14]), .ip2(n22997), .op(n23000) );
  inv_1 U27124 ( .ip(\x[6][14] ), .op(n22998) );
  or2_1 U27125 ( .ip1(n22998), .ip2(n22997), .op(n22999) );
  nand2_1 U27126 ( .ip1(n23000), .ip2(n22999), .op(n23578) );
  nor2_1 U27127 ( .ip1(n23001), .ip2(n23578), .op(n23041) );
  and2_1 U27128 ( .ip1(n24332), .ip2(\x[6][13] ), .op(n23002) );
  not_ab_or_c_or_d U27129 ( .ip1(\x[6][14] ), .ip2(n24327), .ip3(n23002), 
        .ip4(n23001), .op(n23553) );
  nor2_1 U27130 ( .ip1(\x[6][13] ), .ip2(n24376), .op(n23004) );
  nor2_1 U27131 ( .ip1(\x[6][12] ), .ip2(n24450), .op(n23003) );
  nor2_1 U27132 ( .ip1(n23004), .ip2(n23003), .op(n23577) );
  inv_1 U27133 ( .ip(n23577), .op(n23005) );
  nand2_1 U27134 ( .ip1(n23553), .ip2(n23005), .op(n23039) );
  nand2_1 U27135 ( .ip1(\x[6][12] ), .ip2(n24449), .op(n23552) );
  inv_1 U27136 ( .ip(\x[6][11] ), .op(n23034) );
  and2_1 U27137 ( .ip1(n23146), .ip2(\x[6][10] ), .op(n23031) );
  inv_1 U27138 ( .ip(\x[6][9] ), .op(n23029) );
  nor2_1 U27139 ( .ip1(\x[6][8] ), .ip2(n23971), .op(n23028) );
  and2_1 U27140 ( .ip1(n23804), .ip2(\x[6][8] ), .op(n23026) );
  inv_1 U27141 ( .ip(\x[6][6] ), .op(n23024) );
  nor2_1 U27142 ( .ip1(sig_in[6]), .ip2(n23024), .op(n23021) );
  inv_1 U27143 ( .ip(\x[6][3] ), .op(n23014) );
  and2_1 U27144 ( .ip1(n24335), .ip2(\x[6][2] ), .op(n23011) );
  nand2_1 U27145 ( .ip1(\x[6][1] ), .ip2(n20652), .op(n23009) );
  nand2_1 U27146 ( .ip1(\x[6][0] ), .ip2(n24143), .op(n23008) );
  nor2_1 U27147 ( .ip1(\x[6][2] ), .ip2(n24107), .op(n23007) );
  nor2_1 U27148 ( .ip1(\x[6][1] ), .ip2(n20652), .op(n23006) );
  not_ab_or_c_or_d U27149 ( .ip1(n23009), .ip2(n23008), .ip3(n23007), .ip4(
        n23006), .op(n23010) );
  not_ab_or_c_or_d U27150 ( .ip1(\x[6][3] ), .ip2(n22795), .ip3(n23011), .ip4(
        n23010), .op(n23013) );
  nor2_1 U27151 ( .ip1(\x[6][4] ), .ip2(n23860), .op(n23012) );
  not_ab_or_c_or_d U27152 ( .ip1(n23251), .ip2(n23014), .ip3(n23013), .ip4(
        n23012), .op(n23015) );
  or2_1 U27153 ( .ip1(\x[6][4] ), .ip2(n23015), .op(n23017) );
  or2_1 U27154 ( .ip1(n23860), .ip2(n23015), .op(n23016) );
  nand2_1 U27155 ( .ip1(n23017), .ip2(n23016), .op(n23019) );
  nor2_1 U27156 ( .ip1(\x[6][5] ), .ip2(n24350), .op(n23018) );
  nor2_1 U27157 ( .ip1(n23019), .ip2(n23018), .op(n23020) );
  not_ab_or_c_or_d U27158 ( .ip1(\x[6][5] ), .ip2(n24482), .ip3(n23021), .ip4(
        n23020), .op(n23023) );
  nor2_1 U27159 ( .ip1(\x[6][7] ), .ip2(n24492), .op(n23022) );
  not_ab_or_c_or_d U27160 ( .ip1(sig_in[6]), .ip2(n23024), .ip3(n23023), .ip4(
        n23022), .op(n23025) );
  not_ab_or_c_or_d U27161 ( .ip1(\x[6][7] ), .ip2(n24492), .ip3(n23026), .ip4(
        n23025), .op(n23027) );
  not_ab_or_c_or_d U27162 ( .ip1(sig_in[9]), .ip2(n23029), .ip3(n23028), .ip4(
        n23027), .op(n23030) );
  not_ab_or_c_or_d U27163 ( .ip1(\x[6][9] ), .ip2(n24455), .ip3(n23031), .ip4(
        n23030), .op(n23033) );
  nor2_1 U27164 ( .ip1(\x[6][10] ), .ip2(n24370), .op(n23032) );
  not_ab_or_c_or_d U27165 ( .ip1(sig_in[11]), .ip2(n23034), .ip3(n23033), 
        .ip4(n23032), .op(n23035) );
  or2_1 U27166 ( .ip1(\x[6][11] ), .ip2(n23035), .op(n23037) );
  or2_1 U27167 ( .ip1(n24136), .ip2(n23035), .op(n23036) );
  nand2_1 U27168 ( .ip1(n23037), .ip2(n23036), .op(n23575) );
  nand3_1 U27169 ( .ip1(n23553), .ip2(n23552), .ip3(n23575), .op(n23038) );
  nand2_1 U27170 ( .ip1(n23039), .ip2(n23038), .op(n23040) );
  nor4_1 U27171 ( .ip1(n23043), .ip2(n23042), .ip3(n23041), .ip4(n23040), .op(
        n24761) );
  nand2_1 U27172 ( .ip1(\x[8][15] ), .ip2(n24186), .op(n23134) );
  and2_1 U27173 ( .ip1(n23895), .ip2(\x[8][13] ), .op(n23044) );
  nor2_1 U27174 ( .ip1(\x[8][15] ), .ip2(n24090), .op(n23541) );
  not_ab_or_c_or_d U27175 ( .ip1(\x[8][14] ), .ip2(n23938), .ip3(n23044), 
        .ip4(n23541), .op(n23545) );
  nand2_1 U27176 ( .ip1(\x[8][12] ), .ip2(n24450), .op(n23045) );
  nand2_1 U27177 ( .ip1(n23545), .ip2(n23045), .op(n23500) );
  nand2_1 U27178 ( .ip1(\x[8][10] ), .ip2(n23146), .op(n23071) );
  nor2_1 U27179 ( .ip1(\x[8][9] ), .ip2(n24043), .op(n23066) );
  inv_1 U27180 ( .ip(\x[8][8] ), .op(n23046) );
  nor3_1 U27181 ( .ip1(sig_in[8]), .ip2(n23066), .ip3(n23046), .op(n23069) );
  and2_1 U27182 ( .ip1(n24461), .ip2(\x[8][7] ), .op(n23063) );
  inv_1 U27183 ( .ip(\x[8][3] ), .op(n23053) );
  nor2_1 U27184 ( .ip1(\x[8][2] ), .ip2(n23659), .op(n23052) );
  inv_1 U27185 ( .ip(\x[8][1] ), .op(n23048) );
  nor2_1 U27186 ( .ip1(sig_in[1]), .ip2(n23048), .op(n23050) );
  inv_1 U27187 ( .ip(\x[8][0] ), .op(n23047) );
  not_ab_or_c_or_d U27188 ( .ip1(n24467), .ip2(n23048), .ip3(n23195), .ip4(
        n23047), .op(n23049) );
  not_ab_or_c_or_d U27189 ( .ip1(\x[8][2] ), .ip2(n24470), .ip3(n23050), .ip4(
        n23049), .op(n23051) );
  not_ab_or_c_or_d U27190 ( .ip1(n23251), .ip2(n23053), .ip3(n23052), .ip4(
        n23051), .op(n23057) );
  nand2_1 U27191 ( .ip1(\x[8][5] ), .ip2(n24119), .op(n23055) );
  nand2_1 U27192 ( .ip1(\x[8][4] ), .ip2(n23721), .op(n23054) );
  nand2_1 U27193 ( .ip1(n23055), .ip2(n23054), .op(n23056) );
  not_ab_or_c_or_d U27194 ( .ip1(\x[8][3] ), .ip2(n22525), .ip3(n23057), .ip4(
        n23056), .op(n23061) );
  nor2_1 U27195 ( .ip1(\x[8][5] ), .ip2(n24350), .op(n23060) );
  nor2_1 U27196 ( .ip1(\x[8][6] ), .ip2(n24485), .op(n23059) );
  not_ab_or_c_or_d U27197 ( .ip1(\x[8][5] ), .ip2(n23600), .ip3(\x[8][4] ), 
        .ip4(n24256), .op(n23058) );
  nor4_1 U27198 ( .ip1(n23061), .ip2(n23060), .ip3(n23059), .ip4(n23058), .op(
        n23062) );
  not_ab_or_c_or_d U27199 ( .ip1(\x[8][6] ), .ip2(n24485), .ip3(n23063), .ip4(
        n23062), .op(n23067) );
  nor2_1 U27200 ( .ip1(\x[8][7] ), .ip2(n24492), .op(n23065) );
  nor2_1 U27201 ( .ip1(\x[8][8] ), .ip2(n24100), .op(n23064) );
  nor4_1 U27202 ( .ip1(n23067), .ip2(n23066), .ip3(n23065), .ip4(n23064), .op(
        n23068) );
  not_ab_or_c_or_d U27203 ( .ip1(\x[8][9] ), .ip2(n24455), .ip3(n23069), .ip4(
        n23068), .op(n23070) );
  nand2_1 U27204 ( .ip1(n23071), .ip2(n23070), .op(n23077) );
  nor2_1 U27205 ( .ip1(\x[8][10] ), .ip2(n24457), .op(n23072) );
  or2_1 U27206 ( .ip1(sig_in[11]), .ip2(n23072), .op(n23075) );
  inv_1 U27207 ( .ip(\x[8][11] ), .op(n23073) );
  or2_1 U27208 ( .ip1(n23073), .ip2(n23072), .op(n23074) );
  nand2_1 U27209 ( .ip1(n23075), .ip2(n23074), .op(n23076) );
  nand2_1 U27210 ( .ip1(n23077), .ip2(n23076), .op(n23079) );
  nand2_1 U27211 ( .ip1(\x[8][11] ), .ip2(n24371), .op(n23078) );
  nand2_1 U27212 ( .ip1(n23079), .ip2(n23078), .op(n23499) );
  nor2_1 U27213 ( .ip1(\x[8][13] ), .ip2(n24376), .op(n23080) );
  or2_1 U27214 ( .ip1(sig_in[12]), .ip2(n23080), .op(n23083) );
  inv_1 U27215 ( .ip(\x[8][12] ), .op(n23081) );
  or2_1 U27216 ( .ip1(n23081), .ip2(n23080), .op(n23082) );
  nand2_1 U27217 ( .ip1(n23083), .ip2(n23082), .op(n23501) );
  inv_1 U27218 ( .ip(n23134), .op(n23084) );
  or2_1 U27219 ( .ip1(sig_in[14]), .ip2(n23084), .op(n23087) );
  inv_1 U27220 ( .ip(\x[8][14] ), .op(n23085) );
  or2_1 U27221 ( .ip1(n23085), .ip2(n23084), .op(n23086) );
  nand2_1 U27222 ( .ip1(n23087), .ip2(n23086), .op(n23540) );
  and3_1 U27223 ( .ip1(n23499), .ip2(n23501), .ip3(n23540), .op(n23133) );
  nor2_1 U27224 ( .ip1(\x[9][13] ), .ip2(n24081), .op(n23091) );
  nor2_1 U27225 ( .ip1(\x[9][12] ), .ip2(n24233), .op(n23090) );
  nor2_1 U27226 ( .ip1(\x[9][14] ), .ip2(n24327), .op(n23089) );
  and2_1 U27227 ( .ip1(n24186), .ip2(\x[9][15] ), .op(n23088) );
  nor4_1 U27228 ( .ip1(n23091), .ip2(n23090), .ip3(n23089), .ip4(n23088), .op(
        n23489) );
  nor2_1 U27229 ( .ip1(\x[9][15] ), .ip2(n24329), .op(n23487) );
  or2_1 U27230 ( .ip1(n23489), .ip2(n23487), .op(n23131) );
  nand2_1 U27231 ( .ip1(\x[9][11] ), .ip2(n24239), .op(n23129) );
  and2_1 U27232 ( .ip1(n24450), .ip2(\x[9][12] ), .op(n23126) );
  inv_1 U27233 ( .ip(\x[9][9] ), .op(n23117) );
  nor2_1 U27234 ( .ip1(n21171), .ip2(n23117), .op(n23120) );
  and2_1 U27235 ( .ip1(n23804), .ip2(\x[9][8] ), .op(n23114) );
  inv_1 U27236 ( .ip(\x[9][6] ), .op(n23112) );
  inv_1 U27237 ( .ip(\x[9][5] ), .op(n23104) );
  nor2_1 U27238 ( .ip1(sig_in[5]), .ip2(n23104), .op(n23102) );
  inv_1 U27239 ( .ip(\x[9][3] ), .op(n23100) );
  and2_1 U27240 ( .ip1(n24335), .ip2(\x[9][2] ), .op(n23097) );
  nand2_1 U27241 ( .ip1(\x[9][1] ), .ip2(n20652), .op(n23095) );
  nand2_1 U27242 ( .ip1(\x[9][0] ), .ip2(n24143), .op(n23094) );
  nor2_1 U27243 ( .ip1(\x[9][2] ), .ip2(n23659), .op(n23093) );
  nor2_1 U27244 ( .ip1(\x[9][1] ), .ip2(n20652), .op(n23092) );
  not_ab_or_c_or_d U27245 ( .ip1(n23095), .ip2(n23094), .ip3(n23093), .ip4(
        n23092), .op(n23096) );
  not_ab_or_c_or_d U27246 ( .ip1(\x[9][3] ), .ip2(n22795), .ip3(n23097), .ip4(
        n23096), .op(n23099) );
  nor2_1 U27247 ( .ip1(\x[9][4] ), .ip2(n23860), .op(n23098) );
  not_ab_or_c_or_d U27248 ( .ip1(sig_in[3]), .ip2(n23100), .ip3(n23099), .ip4(
        n23098), .op(n23101) );
  not_ab_or_c_or_d U27249 ( .ip1(\x[9][4] ), .ip2(n23860), .ip3(n23102), .ip4(
        n23101), .op(n23103) );
  or2_1 U27250 ( .ip1(sig_in[5]), .ip2(n23103), .op(n23106) );
  or2_1 U27251 ( .ip1(n23104), .ip2(n23103), .op(n23105) );
  nand2_1 U27252 ( .ip1(n23106), .ip2(n23105), .op(n23107) );
  or2_1 U27253 ( .ip1(\x[9][6] ), .ip2(n23107), .op(n23109) );
  or2_1 U27254 ( .ip1(n24355), .ip2(n23107), .op(n23108) );
  nand2_1 U27255 ( .ip1(n23109), .ip2(n23108), .op(n23111) );
  nor2_1 U27256 ( .ip1(\x[9][7] ), .ip2(n24044), .op(n23110) );
  not_ab_or_c_or_d U27257 ( .ip1(sig_in[6]), .ip2(n23112), .ip3(n23111), .ip4(
        n23110), .op(n23113) );
  not_ab_or_c_or_d U27258 ( .ip1(\x[9][7] ), .ip2(n24492), .ip3(n23114), .ip4(
        n23113), .op(n23116) );
  nor2_1 U27259 ( .ip1(\x[9][8] ), .ip2(n23971), .op(n23115) );
  not_ab_or_c_or_d U27260 ( .ip1(sig_in[9]), .ip2(n23117), .ip3(n23116), .ip4(
        n23115), .op(n23119) );
  and2_1 U27261 ( .ip1(n23146), .ip2(\x[9][10] ), .op(n23118) );
  nor3_1 U27262 ( .ip1(n23120), .ip2(n23119), .ip3(n23118), .op(n23124) );
  nor2_1 U27263 ( .ip1(\x[9][11] ), .ip2(n24456), .op(n23122) );
  nor2_1 U27264 ( .ip1(\x[9][10] ), .ip2(n24370), .op(n23121) );
  or2_1 U27265 ( .ip1(n23122), .ip2(n23121), .op(n23123) );
  nor2_1 U27266 ( .ip1(n23124), .ip2(n23123), .op(n23125) );
  not_ab_or_c_or_d U27267 ( .ip1(\x[9][14] ), .ip2(n23938), .ip3(n23126), 
        .ip4(n23125), .op(n23128) );
  nand2_1 U27268 ( .ip1(\x[9][13] ), .ip2(n24235), .op(n23127) );
  nand3_1 U27269 ( .ip1(n23129), .ip2(n23128), .ip3(n23127), .op(n23488) );
  or2_1 U27270 ( .ip1(n23488), .ip2(n23487), .op(n23130) );
  nand2_1 U27271 ( .ip1(n23131), .ip2(n23130), .op(n23132) );
  not_ab_or_c_or_d U27272 ( .ip1(n23134), .ip2(n23500), .ip3(n23133), .ip4(
        n23132), .op(n24742) );
  nand2_1 U27273 ( .ip1(n24329), .ip2(\x[11][15] ), .op(n23453) );
  inv_1 U27274 ( .ip(n23453), .op(n23135) );
  or2_1 U27275 ( .ip1(sig_in[14]), .ip2(n23135), .op(n23138) );
  inv_1 U27276 ( .ip(\x[11][14] ), .op(n23136) );
  or2_1 U27277 ( .ip1(n23136), .ip2(n23135), .op(n23137) );
  nand2_1 U27278 ( .ip1(n23138), .ip2(n23137), .op(n23468) );
  nor2_1 U27279 ( .ip1(\x[11][15] ), .ip2(n24090), .op(n23186) );
  nor2_1 U27280 ( .ip1(n23468), .ip2(n23186), .op(n23227) );
  nand2_1 U27281 ( .ip1(n24230), .ip2(\x[10][14] ), .op(n23140) );
  or2_1 U27282 ( .ip1(n24329), .ip2(\x[10][15] ), .op(n23485) );
  nand2_1 U27283 ( .ip1(\x[10][13] ), .ip2(n24235), .op(n23139) );
  nand3_1 U27284 ( .ip1(n23140), .ip2(n23485), .ip3(n23139), .op(n23494) );
  or2_1 U27285 ( .ip1(\x[10][12] ), .ip2(n23494), .op(n23142) );
  or2_1 U27286 ( .ip1(n24449), .ip2(n23494), .op(n23141) );
  nand2_1 U27287 ( .ip1(n23142), .ip2(n23141), .op(n23145) );
  nand2_1 U27288 ( .ip1(n23143), .ip2(\x[10][15] ), .op(n23179) );
  inv_1 U27289 ( .ip(n23179), .op(n23144) );
  nor2_1 U27290 ( .ip1(n23145), .ip2(n23144), .op(n23226) );
  inv_1 U27291 ( .ip(\x[10][11] ), .op(n23173) );
  and2_1 U27292 ( .ip1(n23146), .ip2(\x[10][10] ), .op(n23170) );
  nor2_1 U27293 ( .ip1(\x[10][7] ), .ip2(n24044), .op(n23161) );
  inv_1 U27294 ( .ip(\x[10][6] ), .op(n23147) );
  nor3_1 U27295 ( .ip1(sig_in[6]), .ip2(n23161), .ip3(n23147), .op(n23164) );
  and2_1 U27296 ( .ip1(n24350), .ip2(\x[10][5] ), .op(n23158) );
  inv_1 U27297 ( .ip(\x[10][3] ), .op(n23156) );
  and2_1 U27298 ( .ip1(n24107), .ip2(\x[10][2] ), .op(n23153) );
  nand2_1 U27299 ( .ip1(\x[10][1] ), .ip2(n21685), .op(n23151) );
  nand2_1 U27300 ( .ip1(\x[10][0] ), .ip2(n24143), .op(n23150) );
  nor2_1 U27301 ( .ip1(\x[10][2] ), .ip2(n23659), .op(n23149) );
  nor2_1 U27302 ( .ip1(\x[10][1] ), .ip2(n21685), .op(n23148) );
  not_ab_or_c_or_d U27303 ( .ip1(n23151), .ip2(n23150), .ip3(n23149), .ip4(
        n23148), .op(n23152) );
  not_ab_or_c_or_d U27304 ( .ip1(\x[10][3] ), .ip2(n24342), .ip3(n23153), 
        .ip4(n23152), .op(n23155) );
  nor2_1 U27305 ( .ip1(\x[10][4] ), .ip2(n24347), .op(n23154) );
  not_ab_or_c_or_d U27306 ( .ip1(n23251), .ip2(n23156), .ip3(n23155), .ip4(
        n23154), .op(n23157) );
  not_ab_or_c_or_d U27307 ( .ip1(\x[10][4] ), .ip2(n23860), .ip3(n23158), 
        .ip4(n23157), .op(n23162) );
  nor2_1 U27308 ( .ip1(\x[10][5] ), .ip2(n24350), .op(n23160) );
  nor2_1 U27309 ( .ip1(\x[10][6] ), .ip2(n24355), .op(n23159) );
  nor4_1 U27310 ( .ip1(n23162), .ip2(n23161), .ip3(n23160), .ip4(n23159), .op(
        n23163) );
  not_ab_or_c_or_d U27311 ( .ip1(\x[10][8] ), .ip2(n24100), .ip3(n23164), 
        .ip4(n23163), .op(n23168) );
  nand2_1 U27312 ( .ip1(\x[10][7] ), .ip2(n24492), .op(n23167) );
  nor2_1 U27313 ( .ip1(\x[10][9] ), .ip2(n24269), .op(n23166) );
  nor2_1 U27314 ( .ip1(\x[10][8] ), .ip2(n23971), .op(n23165) );
  not_ab_or_c_or_d U27315 ( .ip1(n23168), .ip2(n23167), .ip3(n23166), .ip4(
        n23165), .op(n23169) );
  not_ab_or_c_or_d U27316 ( .ip1(\x[10][9] ), .ip2(n23981), .ip3(n23170), 
        .ip4(n23169), .op(n23172) );
  nor2_1 U27317 ( .ip1(\x[10][10] ), .ip2(n23980), .op(n23171) );
  not_ab_or_c_or_d U27318 ( .ip1(sig_in[11]), .ip2(n23173), .ip3(n23172), 
        .ip4(n23171), .op(n23174) );
  or2_1 U27319 ( .ip1(\x[10][11] ), .ip2(n23174), .op(n23176) );
  or2_1 U27320 ( .ip1(n24136), .ip2(n23174), .op(n23175) );
  nand2_1 U27321 ( .ip1(n23176), .ip2(n23175), .op(n23490) );
  nor2_1 U27322 ( .ip1(\x[10][13] ), .ip2(n24137), .op(n23178) );
  nor2_1 U27323 ( .ip1(\x[10][12] ), .ip2(n24449), .op(n23177) );
  nor2_1 U27324 ( .ip1(n23178), .ip2(n23177), .op(n23492) );
  inv_1 U27325 ( .ip(n23492), .op(n23181) );
  or2_1 U27326 ( .ip1(n24382), .ip2(\x[10][14] ), .op(n23180) );
  nand2_1 U27327 ( .ip1(n23180), .ip2(n23179), .op(n23484) );
  nor3_1 U27328 ( .ip1(n23490), .ip2(n23181), .ip3(n23484), .op(n23225) );
  nor2_1 U27329 ( .ip1(\x[11][13] ), .ip2(n24376), .op(n23182) );
  or2_1 U27330 ( .ip1(sig_in[12]), .ip2(n23182), .op(n23185) );
  inv_1 U27331 ( .ip(\x[11][12] ), .op(n23183) );
  or2_1 U27332 ( .ip1(n23183), .ip2(n23182), .op(n23184) );
  nand2_1 U27333 ( .ip1(n23185), .ip2(n23184), .op(n23467) );
  nand2_1 U27334 ( .ip1(n23938), .ip2(\x[11][14] ), .op(n23189) );
  inv_1 U27335 ( .ip(n23186), .op(n23188) );
  nand2_1 U27336 ( .ip1(\x[11][13] ), .ip2(n24235), .op(n23187) );
  nand3_1 U27337 ( .ip1(n23189), .ip2(n23188), .ip3(n23187), .op(n23450) );
  or2_1 U27338 ( .ip1(n23467), .ip2(n23450), .op(n23223) );
  nand2_1 U27339 ( .ip1(\x[11][10] ), .ip2(n23980), .op(n23459) );
  nor2_1 U27340 ( .ip1(\x[11][9] ), .ip2(n23981), .op(n23458) );
  nor2_1 U27341 ( .ip1(\x[11][8] ), .ip2(n24100), .op(n23190) );
  nor2_1 U27342 ( .ip1(n23458), .ip2(n23190), .op(n23466) );
  and2_1 U27343 ( .ip1(\x[11][9] ), .ip2(n24164), .op(n23191) );
  or2_1 U27344 ( .ip1(n23466), .ip2(n23191), .op(n23216) );
  or2_1 U27345 ( .ip1(\x[11][8] ), .ip2(n23191), .op(n23193) );
  or2_1 U27346 ( .ip1(n24491), .ip2(n23191), .op(n23192) );
  nand2_1 U27347 ( .ip1(n23193), .ip2(n23192), .op(n23457) );
  nor2_1 U27348 ( .ip1(n24142), .ip2(\x[11][7] ), .op(n23213) );
  inv_1 U27349 ( .ip(\x[11][3] ), .op(n23201) );
  nor2_1 U27350 ( .ip1(\x[11][2] ), .ip2(n23717), .op(n23200) );
  inv_1 U27351 ( .ip(\x[11][1] ), .op(n23196) );
  nor2_1 U27352 ( .ip1(n24464), .ip2(n23196), .op(n23198) );
  inv_1 U27353 ( .ip(\x[11][0] ), .op(n23194) );
  not_ab_or_c_or_d U27354 ( .ip1(n24464), .ip2(n23196), .ip3(n23195), .ip4(
        n23194), .op(n23197) );
  not_ab_or_c_or_d U27355 ( .ip1(\x[11][2] ), .ip2(n24470), .ip3(n23198), 
        .ip4(n23197), .op(n23199) );
  not_ab_or_c_or_d U27356 ( .ip1(n24251), .ip2(n23201), .ip3(n23200), .ip4(
        n23199), .op(n23205) );
  nand2_1 U27357 ( .ip1(\x[11][5] ), .ip2(n24119), .op(n23203) );
  nand2_1 U27358 ( .ip1(\x[11][4] ), .ip2(n23721), .op(n23202) );
  nand2_1 U27359 ( .ip1(n23203), .ip2(n23202), .op(n23204) );
  not_ab_or_c_or_d U27360 ( .ip1(\x[11][3] ), .ip2(n24342), .ip3(n23205), 
        .ip4(n23204), .op(n23209) );
  nor2_1 U27361 ( .ip1(\x[11][6] ), .ip2(n24355), .op(n23208) );
  nor2_1 U27362 ( .ip1(\x[11][5] ), .ip2(n24350), .op(n23207) );
  not_ab_or_c_or_d U27363 ( .ip1(\x[11][5] ), .ip2(n24482), .ip3(\x[11][4] ), 
        .ip4(n24256), .op(n23206) );
  nor4_1 U27364 ( .ip1(n23209), .ip2(n23208), .ip3(n23207), .ip4(n23206), .op(
        n23211) );
  and2_1 U27365 ( .ip1(n24485), .ip2(\x[11][6] ), .op(n23210) );
  not_ab_or_c_or_d U27366 ( .ip1(\x[11][7] ), .ip2(n24142), .ip3(n23211), 
        .ip4(n23210), .op(n23212) );
  nor2_1 U27367 ( .ip1(n23213), .ip2(n23212), .op(n23465) );
  inv_1 U27368 ( .ip(n23465), .op(n23214) );
  nand2_1 U27369 ( .ip1(n23457), .ip2(n23214), .op(n23215) );
  nand2_1 U27370 ( .ip1(n23216), .ip2(n23215), .op(n23217) );
  nand2_1 U27371 ( .ip1(n23459), .ip2(n23217), .op(n23218) );
  nor2_1 U27372 ( .ip1(\x[11][11] ), .ip2(n24456), .op(n23463) );
  nor2_1 U27373 ( .ip1(\x[11][10] ), .ip2(n23980), .op(n23456) );
  nor2_1 U27374 ( .ip1(n23463), .ip2(n23456), .op(n23464) );
  nand2_1 U27375 ( .ip1(n23218), .ip2(n23464), .op(n23220) );
  nand2_1 U27376 ( .ip1(\x[11][11] ), .ip2(n24371), .op(n23219) );
  nand2_1 U27377 ( .ip1(\x[11][12] ), .ip2(n24450), .op(n23451) );
  nand3_1 U27378 ( .ip1(n23220), .ip2(n23219), .ip3(n23451), .op(n23221) );
  or2_1 U27379 ( .ip1(n23221), .ip2(n23450), .op(n23222) );
  nand2_1 U27380 ( .ip1(n23223), .ip2(n23222), .op(n23224) );
  nor4_1 U27381 ( .ip1(n23227), .ip2(n23226), .ip3(n23225), .ip4(n23224), .op(
        n24745) );
  nand2_1 U27382 ( .ip1(\x[13][15] ), .ip2(n24186), .op(n23322) );
  and2_1 U27383 ( .ip1(n24332), .ip2(\x[13][13] ), .op(n23228) );
  nor2_1 U27384 ( .ip1(\x[13][15] ), .ip2(n24090), .op(n23401) );
  not_ab_or_c_or_d U27385 ( .ip1(\x[13][14] ), .ip2(n24230), .ip3(n23228), 
        .ip4(n23401), .op(n23405) );
  nand2_1 U27386 ( .ip1(\x[13][12] ), .ip2(n24450), .op(n23229) );
  nand2_1 U27387 ( .ip1(n23405), .ip2(n23229), .op(n23398) );
  inv_1 U27388 ( .ip(n23322), .op(n23230) );
  or2_1 U27389 ( .ip1(sig_in[14]), .ip2(n23230), .op(n23233) );
  inv_1 U27390 ( .ip(\x[13][14] ), .op(n23231) );
  or2_1 U27391 ( .ip1(n23231), .ip2(n23230), .op(n23232) );
  nand2_1 U27392 ( .ip1(n23233), .ip2(n23232), .op(n23400) );
  nor2_1 U27393 ( .ip1(\x[13][13] ), .ip2(n24137), .op(n23234) );
  or2_1 U27394 ( .ip1(sig_in[12]), .ip2(n23234), .op(n23237) );
  inv_1 U27395 ( .ip(\x[13][12] ), .op(n23235) );
  or2_1 U27396 ( .ip1(n23235), .ip2(n23234), .op(n23236) );
  nand2_1 U27397 ( .ip1(n23237), .ip2(n23236), .op(n23383) );
  nand2_1 U27398 ( .ip1(\x[13][10] ), .ip2(n23980), .op(n23238) );
  nand2_1 U27399 ( .ip1(\x[13][11] ), .ip2(n24371), .op(n23397) );
  nand2_1 U27400 ( .ip1(n23238), .ip2(n23397), .op(n23390) );
  nor2_1 U27401 ( .ip1(\x[13][9] ), .ip2(n24269), .op(n23242) );
  or2_1 U27402 ( .ip1(sig_in[8]), .ip2(n23242), .op(n23241) );
  inv_1 U27403 ( .ip(\x[13][8] ), .op(n23239) );
  or2_1 U27404 ( .ip1(n23239), .ip2(n23242), .op(n23240) );
  nand2_1 U27405 ( .ip1(n23241), .ip2(n23240), .op(n23393) );
  nand2_1 U27406 ( .ip1(\x[13][9] ), .ip2(n24164), .op(n23389) );
  nand2_1 U27407 ( .ip1(\x[13][8] ), .ip2(n23804), .op(n23388) );
  or2_1 U27408 ( .ip1(n23388), .ip2(n23242), .op(n23243) );
  nand2_1 U27409 ( .ip1(n23389), .ip2(n23243), .op(n23266) );
  or2_1 U27410 ( .ip1(n23393), .ip2(n23266), .op(n23268) );
  inv_1 U27411 ( .ip(\x[13][7] ), .op(n23263) );
  nor2_1 U27412 ( .ip1(sig_in[7]), .ip2(n23263), .op(n23261) );
  inv_1 U27413 ( .ip(\x[13][3] ), .op(n23250) );
  inv_1 U27414 ( .ip(\x[13][1] ), .op(n23245) );
  nor2_1 U27415 ( .ip1(sig_in[1]), .ip2(n23245), .op(n23247) );
  inv_1 U27416 ( .ip(\x[13][0] ), .op(n23244) );
  not_ab_or_c_or_d U27417 ( .ip1(n24464), .ip2(n23245), .ip3(sig_in[0]), .ip4(
        n23244), .op(n23246) );
  not_ab_or_c_or_d U27418 ( .ip1(\x[13][2] ), .ip2(n24470), .ip3(n23247), 
        .ip4(n23246), .op(n23249) );
  nor2_1 U27419 ( .ip1(\x[13][2] ), .ip2(n23717), .op(n23248) );
  not_ab_or_c_or_d U27420 ( .ip1(n23251), .ip2(n23250), .ip3(n23249), .ip4(
        n23248), .op(n23255) );
  nand2_1 U27421 ( .ip1(\x[13][5] ), .ip2(n24119), .op(n23253) );
  nand2_1 U27422 ( .ip1(\x[13][4] ), .ip2(n23721), .op(n23252) );
  nand2_1 U27423 ( .ip1(n23253), .ip2(n23252), .op(n23254) );
  not_ab_or_c_or_d U27424 ( .ip1(\x[13][3] ), .ip2(n22795), .ip3(n23255), 
        .ip4(n23254), .op(n23259) );
  nor2_1 U27425 ( .ip1(\x[13][6] ), .ip2(n24485), .op(n23258) );
  nor2_1 U27426 ( .ip1(\x[13][5] ), .ip2(n24350), .op(n23257) );
  not_ab_or_c_or_d U27427 ( .ip1(\x[13][5] ), .ip2(n23600), .ip3(\x[13][4] ), 
        .ip4(n24256), .op(n23256) );
  nor4_1 U27428 ( .ip1(n23259), .ip2(n23258), .ip3(n23257), .ip4(n23256), .op(
        n23260) );
  not_ab_or_c_or_d U27429 ( .ip1(\x[13][6] ), .ip2(n23509), .ip3(n23261), 
        .ip4(n23260), .op(n23262) );
  or2_1 U27430 ( .ip1(sig_in[7]), .ip2(n23262), .op(n23265) );
  or2_1 U27431 ( .ip1(n23263), .ip2(n23262), .op(n23264) );
  nand2_1 U27432 ( .ip1(n23265), .ip2(n23264), .op(n23386) );
  or2_1 U27433 ( .ip1(n23386), .ip2(n23266), .op(n23267) );
  nand2_1 U27434 ( .ip1(n23268), .ip2(n23267), .op(n23269) );
  nor2_1 U27435 ( .ip1(\x[13][10] ), .ip2(n23980), .op(n23384) );
  nor2_1 U27436 ( .ip1(n23269), .ip2(n23384), .op(n23270) );
  nor2_1 U27437 ( .ip1(n23390), .ip2(n23270), .op(n23271) );
  nor2_1 U27438 ( .ip1(\x[13][11] ), .ip2(n21793), .op(n23385) );
  nor2_1 U27439 ( .ip1(n23271), .ip2(n23385), .op(n23272) );
  and3_1 U27440 ( .ip1(n23400), .ip2(n23383), .ip3(n23272), .op(n23321) );
  nand2_1 U27441 ( .ip1(n24332), .ip2(\x[14][13] ), .op(n23274) );
  nand2_1 U27442 ( .ip1(\x[14][12] ), .ip2(n24450), .op(n23273) );
  nand2_1 U27443 ( .ip1(n23274), .ip2(n23273), .op(n23323) );
  nor2_1 U27444 ( .ip1(n24456), .ip2(\x[14][11] ), .op(n23307) );
  nor2_1 U27445 ( .ip1(\x[14][9] ), .ip2(n24043), .op(n23297) );
  inv_1 U27446 ( .ip(\x[14][8] ), .op(n23299) );
  nor3_1 U27447 ( .ip1(sig_in[8]), .ip2(n23297), .ip3(n23299), .op(n23301) );
  inv_1 U27448 ( .ip(\x[14][6] ), .op(n23293) );
  inv_1 U27449 ( .ip(\x[14][1] ), .op(n23276) );
  inv_1 U27450 ( .ip(\x[14][0] ), .op(n23275) );
  not_ab_or_c_or_d U27451 ( .ip1(n24464), .ip2(n23276), .ip3(sig_in[0]), .ip4(
        n23275), .op(n23278) );
  and2_1 U27452 ( .ip1(n22795), .ip2(\x[14][3] ), .op(n23277) );
  not_ab_or_c_or_d U27453 ( .ip1(\x[14][2] ), .ip2(n24470), .ip3(n23278), 
        .ip4(n23277), .op(n23282) );
  nand2_1 U27454 ( .ip1(\x[14][1] ), .ip2(n21685), .op(n23281) );
  nor2_1 U27455 ( .ip1(\x[14][3] ), .ip2(n24342), .op(n23280) );
  not_ab_or_c_or_d U27456 ( .ip1(\x[14][3] ), .ip2(n24342), .ip3(\x[14][2] ), 
        .ip4(n24107), .op(n23279) );
  not_ab_or_c_or_d U27457 ( .ip1(n23282), .ip2(n23281), .ip3(n23280), .ip4(
        n23279), .op(n23284) );
  nand2_1 U27458 ( .ip1(\x[14][4] ), .ip2(n23284), .op(n23287) );
  nor2_1 U27459 ( .ip1(\x[14][5] ), .ip2(n23283), .op(n23286) );
  nor2_1 U27460 ( .ip1(\x[14][4] ), .ip2(n23284), .op(n23285) );
  ab_or_c_or_d U27461 ( .ip1(sig_in[4]), .ip2(n23287), .ip3(n23286), .ip4(
        n23285), .op(n23290) );
  nand2_1 U27462 ( .ip1(\x[14][6] ), .ip2(n24485), .op(n23289) );
  nand2_1 U27463 ( .ip1(\x[14][5] ), .ip2(n24119), .op(n23288) );
  and3_1 U27464 ( .ip1(n23290), .ip2(n23289), .ip3(n23288), .op(n23292) );
  nor2_1 U27465 ( .ip1(\x[14][7] ), .ip2(n24044), .op(n23291) );
  not_ab_or_c_or_d U27466 ( .ip1(sig_in[6]), .ip2(n23293), .ip3(n23292), .ip4(
        n23291), .op(n23294) );
  or2_1 U27467 ( .ip1(\x[14][7] ), .ip2(n23294), .op(n23296) );
  or2_1 U27468 ( .ip1(n24492), .ip2(n23294), .op(n23295) );
  nand2_1 U27469 ( .ip1(n23296), .ip2(n23295), .op(n23298) );
  not_ab_or_c_or_d U27470 ( .ip1(n23779), .ip2(n23299), .ip3(n23298), .ip4(
        n23297), .op(n23300) );
  not_ab_or_c_or_d U27471 ( .ip1(\x[14][9] ), .ip2(n24455), .ip3(n23301), 
        .ip4(n23300), .op(n23303) );
  nor2_1 U27472 ( .ip1(\x[14][10] ), .ip2(n24457), .op(n23302) );
  nor2_1 U27473 ( .ip1(n23303), .ip2(n23302), .op(n23305) );
  and2_1 U27474 ( .ip1(n24451), .ip2(\x[14][10] ), .op(n23304) );
  not_ab_or_c_or_d U27475 ( .ip1(\x[14][11] ), .ip2(n24136), .ip3(n23305), 
        .ip4(n23304), .op(n23306) );
  nor2_1 U27476 ( .ip1(n23307), .ip2(n23306), .op(n23326) );
  or2_1 U27477 ( .ip1(n23323), .ip2(n23326), .op(n23312) );
  nor2_1 U27478 ( .ip1(\x[14][13] ), .ip2(n24137), .op(n23308) );
  or2_1 U27479 ( .ip1(sig_in[12]), .ip2(n23308), .op(n23311) );
  inv_1 U27480 ( .ip(\x[14][12] ), .op(n23309) );
  or2_1 U27481 ( .ip1(n23309), .ip2(n23308), .op(n23310) );
  nand2_1 U27482 ( .ip1(n23311), .ip2(n23310), .op(n23325) );
  nand2_1 U27483 ( .ip1(n23312), .ip2(n23325), .op(n23314) );
  nor2_1 U27484 ( .ip1(\x[14][15] ), .ip2(n24090), .op(n23380) );
  and2_1 U27485 ( .ip1(n24230), .ip2(\x[14][14] ), .op(n23324) );
  nor2_1 U27486 ( .ip1(n23380), .ip2(n23324), .op(n23313) );
  nand2_1 U27487 ( .ip1(n23314), .ip2(n23313), .op(n23319) );
  nor2_1 U27488 ( .ip1(\x[14][14] ), .ip2(n23938), .op(n23315) );
  or2_1 U27489 ( .ip1(\x[14][15] ), .ip2(n23315), .op(n23317) );
  or2_1 U27490 ( .ip1(n24384), .ip2(n23315), .op(n23316) );
  nand2_1 U27491 ( .ip1(n23317), .ip2(n23316), .op(n23327) );
  or2_1 U27492 ( .ip1(n23380), .ip2(n23327), .op(n23318) );
  nand2_1 U27493 ( .ip1(n23319), .ip2(n23318), .op(n23320) );
  not_ab_or_c_or_d U27494 ( .ip1(n23322), .ip2(n23398), .ip3(n23321), .ip4(
        n23320), .op(n27420) );
  not_ab_or_c_or_d U27495 ( .ip1(n23326), .ip2(n23325), .ip3(n23324), .ip4(
        n23323), .op(n23329) );
  inv_1 U27496 ( .ip(n23327), .op(n23328) );
  nor2_1 U27497 ( .ip1(n23329), .ip2(n23328), .op(n23379) );
  nor2_1 U27498 ( .ip1(\x[15][15] ), .ip2(n24090), .op(n23372) );
  nand2_1 U27499 ( .ip1(n24384), .ip2(\x[15][15] ), .op(n23710) );
  inv_1 U27500 ( .ip(n23710), .op(n23330) );
  or2_1 U27501 ( .ip1(sig_in[14]), .ip2(n23330), .op(n23333) );
  inv_1 U27502 ( .ip(\x[15][14] ), .op(n23331) );
  or2_1 U27503 ( .ip1(n23331), .ip2(n23330), .op(n23332) );
  nand2_1 U27504 ( .ip1(n23333), .ip2(n23332), .op(n23653) );
  nor2_1 U27505 ( .ip1(n23372), .ip2(n23653), .op(n23378) );
  nor2_1 U27506 ( .ip1(\x[15][13] ), .ip2(n24137), .op(n23335) );
  nor2_1 U27507 ( .ip1(\x[15][12] ), .ip2(n24450), .op(n23334) );
  nor2_1 U27508 ( .ip1(n23335), .ip2(n23334), .op(n23654) );
  inv_1 U27509 ( .ip(n23654), .op(n23371) );
  and2_1 U27510 ( .ip1(n24079), .ip2(\x[15][12] ), .op(n23651) );
  nand2_1 U27511 ( .ip1(\x[15][10] ), .ip2(n24370), .op(n23361) );
  nor2_1 U27512 ( .ip1(\x[15][9] ), .ip2(n24164), .op(n23356) );
  inv_1 U27513 ( .ip(\x[15][8] ), .op(n23336) );
  nor3_1 U27514 ( .ip1(sig_in[8]), .ip2(n23356), .ip3(n23336), .op(n23359) );
  and2_1 U27515 ( .ip1(n24461), .ip2(\x[15][7] ), .op(n23353) );
  inv_1 U27516 ( .ip(\x[15][3] ), .op(n23343) );
  inv_1 U27517 ( .ip(\x[15][1] ), .op(n23338) );
  nor2_1 U27518 ( .ip1(n24464), .ip2(n23338), .op(n23340) );
  inv_1 U27519 ( .ip(\x[15][0] ), .op(n23337) );
  not_ab_or_c_or_d U27520 ( .ip1(n24464), .ip2(n23338), .ip3(sig_in[0]), .ip4(
        n23337), .op(n23339) );
  not_ab_or_c_or_d U27521 ( .ip1(\x[15][2] ), .ip2(n24470), .ip3(n23340), 
        .ip4(n23339), .op(n23342) );
  nor2_1 U27522 ( .ip1(\x[15][2] ), .ip2(n23717), .op(n23341) );
  not_ab_or_c_or_d U27523 ( .ip1(n23251), .ip2(n23343), .ip3(n23342), .ip4(
        n23341), .op(n23347) );
  nand2_1 U27524 ( .ip1(\x[15][5] ), .ip2(n24119), .op(n23345) );
  nand2_1 U27525 ( .ip1(\x[15][4] ), .ip2(n23860), .op(n23344) );
  nand2_1 U27526 ( .ip1(n23345), .ip2(n23344), .op(n23346) );
  not_ab_or_c_or_d U27527 ( .ip1(\x[15][3] ), .ip2(n24476), .ip3(n23347), 
        .ip4(n23346), .op(n23351) );
  nor2_1 U27528 ( .ip1(\x[15][6] ), .ip2(n24355), .op(n23350) );
  nor2_1 U27529 ( .ip1(\x[15][5] ), .ip2(n24350), .op(n23349) );
  not_ab_or_c_or_d U27530 ( .ip1(\x[15][5] ), .ip2(n24482), .ip3(\x[15][4] ), 
        .ip4(n24256), .op(n23348) );
  nor4_1 U27531 ( .ip1(n23351), .ip2(n23350), .ip3(n23349), .ip4(n23348), .op(
        n23352) );
  not_ab_or_c_or_d U27532 ( .ip1(\x[15][6] ), .ip2(n24485), .ip3(n23353), 
        .ip4(n23352), .op(n23357) );
  nor2_1 U27533 ( .ip1(\x[15][7] ), .ip2(n24492), .op(n23355) );
  nor2_1 U27534 ( .ip1(\x[15][8] ), .ip2(n23971), .op(n23354) );
  nor4_1 U27535 ( .ip1(n23357), .ip2(n23356), .ip3(n23355), .ip4(n23354), .op(
        n23358) );
  not_ab_or_c_or_d U27536 ( .ip1(\x[15][9] ), .ip2(n24164), .ip3(n23359), 
        .ip4(n23358), .op(n23360) );
  nand2_1 U27537 ( .ip1(n23361), .ip2(n23360), .op(n23367) );
  nor2_1 U27538 ( .ip1(\x[15][10] ), .ip2(n23980), .op(n23362) );
  or2_1 U27539 ( .ip1(sig_in[11]), .ip2(n23362), .op(n23365) );
  inv_1 U27540 ( .ip(\x[15][11] ), .op(n23363) );
  or2_1 U27541 ( .ip1(n23363), .ip2(n23362), .op(n23364) );
  nand2_1 U27542 ( .ip1(n23365), .ip2(n23364), .op(n23366) );
  nand2_1 U27543 ( .ip1(n23367), .ip2(n23366), .op(n23369) );
  nand2_1 U27544 ( .ip1(\x[15][11] ), .ip2(n24239), .op(n23368) );
  nand2_1 U27545 ( .ip1(n23369), .ip2(n23368), .op(n23655) );
  nor2_1 U27546 ( .ip1(n23651), .ip2(n23655), .op(n23370) );
  nor2_1 U27547 ( .ip1(n23371), .ip2(n23370), .op(n23376) );
  nand2_1 U27548 ( .ip1(n24327), .ip2(\x[15][14] ), .op(n23375) );
  inv_1 U27549 ( .ip(n23372), .op(n23374) );
  nand2_1 U27550 ( .ip1(\x[15][13] ), .ip2(n24081), .op(n23373) );
  nand3_1 U27551 ( .ip1(n23375), .ip2(n23374), .ip3(n23373), .op(n23652) );
  nor2_1 U27552 ( .ip1(n23376), .ip2(n23652), .op(n23377) );
  nor4_1 U27553 ( .ip1(n23380), .ip2(n23379), .ip3(n23378), .ip4(n23377), .op(
        n27419) );
  nor2_1 U27554 ( .ip1(n27420), .ip2(n27419), .op(n24736) );
  and2_1 U27555 ( .ip1(n23895), .ip2(\x[12][13] ), .op(n23381) );
  nor2_1 U27556 ( .ip1(\x[12][15] ), .ip2(n24090), .op(n23474) );
  not_ab_or_c_or_d U27557 ( .ip1(\x[12][14] ), .ip2(n24230), .ip3(n23381), 
        .ip4(n23474), .op(n23478) );
  nand2_1 U27558 ( .ip1(\x[12][12] ), .ip2(n24450), .op(n23382) );
  nand2_1 U27559 ( .ip1(n23478), .ip2(n23382), .op(n23480) );
  nand2_1 U27560 ( .ip1(\x[12][15] ), .ip2(n24186), .op(n23406) );
  nand2_1 U27561 ( .ip1(n23480), .ip2(n23406), .op(n23449) );
  inv_1 U27562 ( .ip(n23383), .op(n23404) );
  or2_1 U27563 ( .ip1(n23385), .ip2(n23384), .op(n23395) );
  inv_1 U27564 ( .ip(n23386), .op(n23387) );
  nand2_1 U27565 ( .ip1(n23388), .ip2(n23387), .op(n23392) );
  inv_1 U27566 ( .ip(n23389), .op(n23391) );
  not_ab_or_c_or_d U27567 ( .ip1(n23393), .ip2(n23392), .ip3(n23391), .ip4(
        n23390), .op(n23394) );
  or2_1 U27568 ( .ip1(n23395), .ip2(n23394), .op(n23396) );
  nand2_1 U27569 ( .ip1(n23397), .ip2(n23396), .op(n23399) );
  nor2_1 U27570 ( .ip1(n23399), .ip2(n23398), .op(n23403) );
  nor2_1 U27571 ( .ip1(n23401), .ip2(n23400), .op(n23402) );
  not_ab_or_c_or_d U27572 ( .ip1(n23405), .ip2(n23404), .ip3(n23403), .ip4(
        n23402), .op(n23448) );
  inv_1 U27573 ( .ip(n23406), .op(n23407) );
  or2_1 U27574 ( .ip1(sig_in[14]), .ip2(n23407), .op(n23410) );
  inv_1 U27575 ( .ip(\x[12][14] ), .op(n23408) );
  or2_1 U27576 ( .ip1(n23408), .ip2(n23407), .op(n23409) );
  nand2_1 U27577 ( .ip1(n23410), .ip2(n23409), .op(n23473) );
  nor2_1 U27578 ( .ip1(\x[12][13] ), .ip2(n24137), .op(n23411) );
  or2_1 U27579 ( .ip1(sig_in[12]), .ip2(n23411), .op(n23414) );
  inv_1 U27580 ( .ip(\x[12][12] ), .op(n23412) );
  or2_1 U27581 ( .ip1(n23412), .ip2(n23411), .op(n23413) );
  nand2_1 U27582 ( .ip1(n23414), .ip2(n23413), .op(n23455) );
  inv_1 U27583 ( .ip(\x[12][11] ), .op(n23444) );
  nor2_1 U27584 ( .ip1(n23444), .ip2(n17981), .op(n23446) );
  and2_1 U27585 ( .ip1(n24451), .ip2(\x[12][10] ), .op(n23441) );
  inv_1 U27586 ( .ip(\x[12][9] ), .op(n23439) );
  nor2_1 U27587 ( .ip1(\x[12][8] ), .ip2(n24100), .op(n23438) );
  nand2_1 U27588 ( .ip1(\x[12][7] ), .ip2(n24461), .op(n23417) );
  nand2_1 U27589 ( .ip1(\x[12][6] ), .ip2(n23770), .op(n23415) );
  nor2_1 U27590 ( .ip1(\x[12][7] ), .ip2(n24044), .op(n23433) );
  or2_1 U27591 ( .ip1(n23415), .ip2(n23433), .op(n23416) );
  nand2_1 U27592 ( .ip1(n23417), .ip2(n23416), .op(n23436) );
  nor2_1 U27593 ( .ip1(\x[12][6] ), .ip2(n24355), .op(n23434) );
  nor2_1 U27594 ( .ip1(\x[12][5] ), .ip2(n24350), .op(n23432) );
  and2_1 U27595 ( .ip1(n24256), .ip2(\x[12][4] ), .op(n23426) );
  inv_1 U27596 ( .ip(\x[12][3] ), .op(n23424) );
  nor2_1 U27597 ( .ip1(\x[12][2] ), .ip2(n23717), .op(n23423) );
  inv_1 U27598 ( .ip(\x[12][1] ), .op(n23419) );
  nor2_1 U27599 ( .ip1(sig_in[1]), .ip2(n23419), .op(n23421) );
  inv_1 U27600 ( .ip(\x[12][0] ), .op(n23418) );
  not_ab_or_c_or_d U27601 ( .ip1(sig_in[1]), .ip2(n23419), .ip3(sig_in[0]), 
        .ip4(n23418), .op(n23420) );
  not_ab_or_c_or_d U27602 ( .ip1(\x[12][2] ), .ip2(n24470), .ip3(n23421), 
        .ip4(n23420), .op(n23422) );
  not_ab_or_c_or_d U27603 ( .ip1(sig_in[3]), .ip2(n23424), .ip3(n23423), .ip4(
        n23422), .op(n23425) );
  not_ab_or_c_or_d U27604 ( .ip1(\x[12][3] ), .ip2(n22795), .ip3(n23426), 
        .ip4(n23425), .op(n23428) );
  nor2_1 U27605 ( .ip1(n24347), .ip2(\x[12][4] ), .op(n23427) );
  nor2_1 U27606 ( .ip1(n23428), .ip2(n23427), .op(n23430) );
  and2_1 U27607 ( .ip1(n23283), .ip2(\x[12][5] ), .op(n23429) );
  nor2_1 U27608 ( .ip1(n23430), .ip2(n23429), .op(n23431) );
  nor4_1 U27609 ( .ip1(n23434), .ip2(n23433), .ip3(n23432), .ip4(n23431), .op(
        n23435) );
  not_ab_or_c_or_d U27610 ( .ip1(\x[12][8] ), .ip2(n24491), .ip3(n23436), 
        .ip4(n23435), .op(n23437) );
  not_ab_or_c_or_d U27611 ( .ip1(sig_in[9]), .ip2(n23439), .ip3(n23438), .ip4(
        n23437), .op(n23440) );
  not_ab_or_c_or_d U27612 ( .ip1(\x[12][9] ), .ip2(n24043), .ip3(n23441), 
        .ip4(n23440), .op(n23443) );
  nor2_1 U27613 ( .ip1(\x[12][10] ), .ip2(n23980), .op(n23442) );
  not_ab_or_c_or_d U27614 ( .ip1(sig_in[11]), .ip2(n23444), .ip3(n23443), 
        .ip4(n23442), .op(n23445) );
  or2_1 U27615 ( .ip1(n23446), .ip2(n23445), .op(n23479) );
  nand3_1 U27616 ( .ip1(n23473), .ip2(n23455), .ip3(n23479), .op(n23447) );
  nand3_1 U27617 ( .ip1(n23449), .ip2(n23448), .ip3(n23447), .op(n24737) );
  inv_1 U27618 ( .ip(n23450), .op(n23452) );
  nand2_1 U27619 ( .ip1(n23452), .ip2(n23451), .op(n23454) );
  nand2_1 U27620 ( .ip1(n23454), .ip2(n23453), .op(n23483) );
  inv_1 U27621 ( .ip(n23455), .op(n23477) );
  nor3_1 U27622 ( .ip1(n23458), .ip2(n23457), .ip3(n23456), .op(n23461) );
  inv_1 U27623 ( .ip(n23459), .op(n23460) );
  not_ab_or_c_or_d U27624 ( .ip1(\x[11][11] ), .ip2(n24136), .ip3(n23461), 
        .ip4(n23460), .op(n23462) );
  or2_1 U27625 ( .ip1(n23463), .ip2(n23462), .op(n23472) );
  nand3_1 U27626 ( .ip1(n23466), .ip2(n23465), .ip3(n23464), .op(n23471) );
  inv_1 U27627 ( .ip(n23467), .op(n23470) );
  inv_1 U27628 ( .ip(n23468), .op(n23469) );
  not_ab_or_c_or_d U27629 ( .ip1(n23472), .ip2(n23471), .ip3(n23470), .ip4(
        n23469), .op(n23476) );
  nor2_1 U27630 ( .ip1(n23474), .ip2(n23473), .op(n23475) );
  not_ab_or_c_or_d U27631 ( .ip1(n23478), .ip2(n23477), .ip3(n23476), .ip4(
        n23475), .op(n23482) );
  or2_1 U27632 ( .ip1(n23480), .ip2(n23479), .op(n23481) );
  nand3_1 U27633 ( .ip1(n23483), .ip2(n23482), .ip3(n23481), .op(n24748) );
  nand3_1 U27634 ( .ip1(n24736), .ip2(n24737), .ip3(n24748), .op(n24746) );
  nor2_1 U27635 ( .ip1(n24745), .ip2(n24746), .op(n24731) );
  and2_1 U27636 ( .ip1(n23485), .ip2(n23484), .op(n23486) );
  not_ab_or_c_or_d U27637 ( .ip1(n23489), .ip2(n23488), .ip3(n23487), .ip4(
        n23486), .op(n23498) );
  nand2_1 U27638 ( .ip1(\x[10][12] ), .ip2(n24450), .op(n23491) );
  nand2_1 U27639 ( .ip1(n23491), .ip2(n23490), .op(n23493) );
  nand2_1 U27640 ( .ip1(n23493), .ip2(n23492), .op(n23496) );
  inv_1 U27641 ( .ip(n23494), .op(n23495) );
  nand2_1 U27642 ( .ip1(n23496), .ip2(n23495), .op(n23497) );
  nand2_1 U27643 ( .ip1(n23498), .ip2(n23497), .op(n24733) );
  nand2_1 U27644 ( .ip1(n24731), .ip2(n24733), .op(n24743) );
  nor2_1 U27645 ( .ip1(n24742), .ip2(n24743), .op(n24734) );
  or2_1 U27646 ( .ip1(n23500), .ip2(n23499), .op(n23551) );
  inv_1 U27647 ( .ip(n23501), .op(n23544) );
  and2_1 U27648 ( .ip1(n24451), .ip2(\x[7][10] ), .op(n23502) );
  and2_1 U27649 ( .ip1(n24239), .ip2(\x[7][11] ), .op(n23506) );
  not_ab_or_c_or_d U27650 ( .ip1(\x[7][9] ), .ip2(n24269), .ip3(n23502), .ip4(
        n23506), .op(n23559) );
  inv_1 U27651 ( .ip(\x[7][8] ), .op(n23531) );
  nor2_1 U27652 ( .ip1(n24455), .ip2(\x[7][9] ), .op(n23530) );
  or3_1 U27653 ( .ip1(n23779), .ip2(n23531), .ip3(n23530), .op(n23503) );
  nand2_1 U27654 ( .ip1(n23559), .ip2(n23503), .op(n23508) );
  nor2_1 U27655 ( .ip1(\x[7][11] ), .ip2(n24456), .op(n23505) );
  nor2_1 U27656 ( .ip1(\x[7][10] ), .ip2(n24370), .op(n23504) );
  nor2_1 U27657 ( .ip1(n23505), .ip2(n23504), .op(n23534) );
  nor2_1 U27658 ( .ip1(n23506), .ip2(n23534), .op(n23566) );
  inv_1 U27659 ( .ip(n23566), .op(n23507) );
  nand2_1 U27660 ( .ip1(n23508), .ip2(n23507), .op(n23539) );
  and2_1 U27661 ( .ip1(n24461), .ip2(\x[7][7] ), .op(n23527) );
  nor2_1 U27662 ( .ip1(n23509), .ip2(\x[7][6] ), .op(n23525) );
  and2_1 U27663 ( .ip1(n24119), .ip2(\x[7][5] ), .op(n23523) );
  nor2_1 U27664 ( .ip1(\x[7][4] ), .ip2(n23721), .op(n23521) );
  and2_1 U27665 ( .ip1(n23860), .ip2(\x[7][4] ), .op(n23518) );
  inv_1 U27666 ( .ip(\x[7][3] ), .op(n23516) );
  nor2_1 U27667 ( .ip1(\x[7][2] ), .ip2(n24107), .op(n23515) );
  inv_1 U27668 ( .ip(\x[7][1] ), .op(n23511) );
  nor2_1 U27669 ( .ip1(n24464), .ip2(n23511), .op(n23513) );
  inv_1 U27670 ( .ip(\x[7][0] ), .op(n23510) );
  not_ab_or_c_or_d U27671 ( .ip1(n24464), .ip2(n23511), .ip3(sig_in[0]), .ip4(
        n23510), .op(n23512) );
  not_ab_or_c_or_d U27672 ( .ip1(\x[7][2] ), .ip2(n24470), .ip3(n23513), .ip4(
        n23512), .op(n23514) );
  not_ab_or_c_or_d U27673 ( .ip1(n24251), .ip2(n23516), .ip3(n23515), .ip4(
        n23514), .op(n23517) );
  not_ab_or_c_or_d U27674 ( .ip1(\x[7][3] ), .ip2(n24342), .ip3(n23518), .ip4(
        n23517), .op(n23520) );
  nor2_1 U27675 ( .ip1(\x[7][5] ), .ip2(n24350), .op(n23519) );
  nor3_1 U27676 ( .ip1(n23521), .ip2(n23520), .ip3(n23519), .op(n23522) );
  nor2_1 U27677 ( .ip1(n23523), .ip2(n23522), .op(n23524) );
  nor2_1 U27678 ( .ip1(n23525), .ip2(n23524), .op(n23526) );
  not_ab_or_c_or_d U27679 ( .ip1(\x[7][6] ), .ip2(n24485), .ip3(n23527), .ip4(
        n23526), .op(n23529) );
  nor2_1 U27680 ( .ip1(\x[7][7] ), .ip2(n24044), .op(n23528) );
  nor2_1 U27681 ( .ip1(n23529), .ip2(n23528), .op(n23562) );
  or2_1 U27682 ( .ip1(sig_in[8]), .ip2(n23530), .op(n23533) );
  or2_1 U27683 ( .ip1(n23531), .ip2(n23530), .op(n23532) );
  nand2_1 U27684 ( .ip1(n23533), .ip2(n23532), .op(n23564) );
  nand3_1 U27685 ( .ip1(n23534), .ip2(n23562), .ip3(n23564), .op(n23538) );
  nor2_1 U27686 ( .ip1(\x[7][13] ), .ip2(n24376), .op(n23536) );
  nor2_1 U27687 ( .ip1(\x[7][12] ), .ip2(n24449), .op(n23535) );
  or2_1 U27688 ( .ip1(n23536), .ip2(n23535), .op(n23573) );
  nand2_1 U27689 ( .ip1(\x[7][15] ), .ip2(n24186), .op(n23548) );
  or2_1 U27690 ( .ip1(n24185), .ip2(\x[7][14] ), .op(n23537) );
  nand2_1 U27691 ( .ip1(n23548), .ip2(n23537), .op(n23556) );
  not_ab_or_c_or_d U27692 ( .ip1(n23539), .ip2(n23538), .ip3(n23573), .ip4(
        n23556), .op(n23543) );
  nor2_1 U27693 ( .ip1(n23541), .ip2(n23540), .op(n23542) );
  not_ab_or_c_or_d U27694 ( .ip1(n23545), .ip2(n23544), .ip3(n23543), .ip4(
        n23542), .op(n23550) );
  and2_1 U27695 ( .ip1(n24332), .ip2(\x[7][13] ), .op(n23546) );
  nor2_1 U27696 ( .ip1(\x[7][15] ), .ip2(n24090), .op(n23557) );
  not_ab_or_c_or_d U27697 ( .ip1(\x[7][14] ), .ip2(n23938), .ip3(n23546), 
        .ip4(n23557), .op(n23574) );
  nand2_1 U27698 ( .ip1(\x[7][12] ), .ip2(n24079), .op(n23547) );
  nand2_1 U27699 ( .ip1(n23574), .ip2(n23547), .op(n23569) );
  nand2_1 U27700 ( .ip1(n23548), .ip2(n23569), .op(n23549) );
  nand3_1 U27701 ( .ip1(n23551), .ip2(n23550), .ip3(n23549), .op(n24735) );
  nand2_1 U27702 ( .ip1(n23553), .ip2(n23552), .op(n23555) );
  nand2_1 U27703 ( .ip1(n23555), .ip2(n23554), .op(n23581) );
  inv_1 U27704 ( .ip(n23556), .op(n23558) );
  nor2_1 U27705 ( .ip1(n23558), .ip2(n23557), .op(n23572) );
  inv_1 U27706 ( .ip(n23559), .op(n23563) );
  or2_1 U27707 ( .ip1(\x[7][8] ), .ip2(n23563), .op(n23561) );
  or2_1 U27708 ( .ip1(n24491), .ip2(n23563), .op(n23560) );
  nand2_1 U27709 ( .ip1(n23561), .ip2(n23560), .op(n23568) );
  inv_1 U27710 ( .ip(n23562), .op(n23567) );
  nor2_1 U27711 ( .ip1(n23564), .ip2(n23563), .op(n23565) );
  not_ab_or_c_or_d U27712 ( .ip1(n23568), .ip2(n23567), .ip3(n23566), .ip4(
        n23565), .op(n23570) );
  nor2_1 U27713 ( .ip1(n23570), .ip2(n23569), .op(n23571) );
  not_ab_or_c_or_d U27714 ( .ip1(n23574), .ip2(n23573), .ip3(n23572), .ip4(
        n23571), .op(n23580) );
  inv_1 U27715 ( .ip(n23575), .op(n23576) );
  nand3_1 U27716 ( .ip1(n23578), .ip2(n23577), .ip3(n23576), .op(n23579) );
  nand3_1 U27717 ( .ip1(n23581), .ip2(n23580), .ip3(n23579), .op(n24750) );
  nand3_1 U27718 ( .ip1(n24734), .ip2(n24735), .ip3(n24750), .op(n24765) );
  nor3_1 U27719 ( .ip1(n24763), .ip2(n24761), .ip3(n24765), .op(n24725) );
  nand2_1 U27720 ( .ip1(n24327), .ip2(\x[3][14] ), .op(n23584) );
  nor2_1 U27721 ( .ip1(n24384), .ip2(\x[3][15] ), .op(n23632) );
  inv_1 U27722 ( .ip(n23632), .op(n23583) );
  nand2_1 U27723 ( .ip1(\x[3][13] ), .ip2(n24235), .op(n23582) );
  nand3_1 U27724 ( .ip1(n23584), .ip2(n23583), .ip3(n23582), .op(n23618) );
  nor2_1 U27725 ( .ip1(\x[3][13] ), .ip2(n24376), .op(n23586) );
  nor2_1 U27726 ( .ip1(\x[3][12] ), .ip2(n24449), .op(n23585) );
  nor2_1 U27727 ( .ip1(n23586), .ip2(n23585), .op(n23646) );
  or2_1 U27728 ( .ip1(n23618), .ip2(n23646), .op(n23634) );
  nand2_1 U27729 ( .ip1(\x[3][11] ), .ip2(n24239), .op(n23615) );
  nand2_1 U27730 ( .ip1(\x[3][10] ), .ip2(n24370), .op(n23614) );
  nor2_1 U27731 ( .ip1(\x[3][5] ), .ip2(n23283), .op(n23596) );
  inv_1 U27732 ( .ip(\x[3][4] ), .op(n23587) );
  nor3_1 U27733 ( .ip1(sig_in[4]), .ip2(n23596), .ip3(n23587), .op(n23599) );
  and2_1 U27734 ( .ip1(n24335), .ip2(\x[3][2] ), .op(n23593) );
  nand2_1 U27735 ( .ip1(\x[3][1] ), .ip2(n21685), .op(n23591) );
  nand2_1 U27736 ( .ip1(\x[3][0] ), .ip2(n24143), .op(n23590) );
  nor2_1 U27737 ( .ip1(\x[3][2] ), .ip2(n23717), .op(n23589) );
  nor2_1 U27738 ( .ip1(\x[3][1] ), .ip2(n20652), .op(n23588) );
  not_ab_or_c_or_d U27739 ( .ip1(n23591), .ip2(n23590), .ip3(n23589), .ip4(
        n23588), .op(n23592) );
  not_ab_or_c_or_d U27740 ( .ip1(\x[3][3] ), .ip2(n24342), .ip3(n23593), .ip4(
        n23592), .op(n23597) );
  nor2_1 U27741 ( .ip1(\x[3][4] ), .ip2(n24256), .op(n23595) );
  nor2_1 U27742 ( .ip1(\x[3][3] ), .ip2(n24476), .op(n23594) );
  nor4_1 U27743 ( .ip1(n23597), .ip2(n23596), .ip3(n23595), .ip4(n23594), .op(
        n23598) );
  not_ab_or_c_or_d U27744 ( .ip1(\x[3][5] ), .ip2(n23600), .ip3(n23599), .ip4(
        n23598), .op(n23604) );
  nand2_1 U27745 ( .ip1(\x[3][6] ), .ip2(n24485), .op(n23603) );
  nor2_1 U27746 ( .ip1(\x[3][6] ), .ip2(n24355), .op(n23602) );
  nor2_1 U27747 ( .ip1(\x[3][7] ), .ip2(n24492), .op(n23601) );
  not_ab_or_c_or_d U27748 ( .ip1(n23604), .ip2(n23603), .ip3(n23602), .ip4(
        n23601), .op(n23608) );
  nand2_1 U27749 ( .ip1(\x[3][9] ), .ip2(n24455), .op(n23606) );
  nand2_1 U27750 ( .ip1(\x[3][8] ), .ip2(n24100), .op(n23605) );
  nand2_1 U27751 ( .ip1(n23606), .ip2(n23605), .op(n23607) );
  not_ab_or_c_or_d U27752 ( .ip1(\x[3][7] ), .ip2(n24492), .ip3(n23608), .ip4(
        n23607), .op(n23612) );
  not_ab_or_c_or_d U27753 ( .ip1(\x[3][9] ), .ip2(n24455), .ip3(\x[3][8] ), 
        .ip4(n24358), .op(n23611) );
  nor2_1 U27754 ( .ip1(\x[3][9] ), .ip2(n24164), .op(n23610) );
  nor2_1 U27755 ( .ip1(\x[3][10] ), .ip2(n24457), .op(n23609) );
  or4_1 U27756 ( .ip1(n23612), .ip2(n23611), .ip3(n23610), .ip4(n23609), .op(
        n23613) );
  nand3_1 U27757 ( .ip1(n23615), .ip2(n23614), .ip3(n23613), .op(n23617) );
  or2_1 U27758 ( .ip1(n24136), .ip2(\x[3][11] ), .op(n23616) );
  nand2_1 U27759 ( .ip1(n23617), .ip2(n23616), .op(n23645) );
  or2_1 U27760 ( .ip1(\x[3][12] ), .ip2(n23618), .op(n23620) );
  or2_1 U27761 ( .ip1(n24449), .ip2(n23618), .op(n23619) );
  nand2_1 U27762 ( .ip1(n23620), .ip2(n23619), .op(n23635) );
  nor2_1 U27763 ( .ip1(n23622), .ip2(n23621), .op(n23623) );
  nor2_1 U27764 ( .ip1(n23624), .ip2(n23623), .op(n23628) );
  nor2_1 U27765 ( .ip1(n23626), .ip2(n23625), .op(n23627) );
  not_ab_or_c_or_d U27766 ( .ip1(n23645), .ip2(n23635), .ip3(n23628), .ip4(
        n23627), .op(n23633) );
  nor2_1 U27767 ( .ip1(\x[3][14] ), .ip2(n23938), .op(n23629) );
  or2_1 U27768 ( .ip1(\x[3][15] ), .ip2(n23629), .op(n23631) );
  or2_1 U27769 ( .ip1(n24329), .ip2(n23629), .op(n23630) );
  nand2_1 U27770 ( .ip1(n23631), .ip2(n23630), .op(n23647) );
  or2_1 U27771 ( .ip1(n23632), .ip2(n23647), .op(n23643) );
  nand3_1 U27772 ( .ip1(n23634), .ip2(n23633), .ip3(n23643), .op(n24726) );
  inv_1 U27773 ( .ip(n23635), .op(n23644) );
  inv_1 U27774 ( .ip(n23636), .op(n23637) );
  nor2_1 U27775 ( .ip1(n23638), .ip2(n23637), .op(n23642) );
  nor2_1 U27776 ( .ip1(n23640), .ip2(n23639), .op(n23641) );
  not_ab_or_c_or_d U27777 ( .ip1(n23644), .ip2(n23643), .ip3(n23642), .ip4(
        n23641), .op(n23650) );
  inv_1 U27778 ( .ip(n23645), .op(n23648) );
  nand3_1 U27779 ( .ip1(n23648), .ip2(n23647), .ip3(n23646), .op(n23649) );
  nand2_1 U27780 ( .ip1(n23650), .ip2(n23649), .op(n24727) );
  nand3_1 U27781 ( .ip1(n24725), .ip2(n24726), .ip3(n24727), .op(n24760) );
  nor2_1 U27782 ( .ip1(n24758), .ip2(n24760), .op(n27436) );
  or2_1 U27783 ( .ip1(n23652), .ip2(n23651), .op(n23711) );
  and3_1 U27784 ( .ip1(n23655), .ip2(n23654), .ip3(n23653), .op(n23709) );
  and2_1 U27785 ( .ip1(n23895), .ip2(\x[16][13] ), .op(n23656) );
  or2_1 U27786 ( .ip1(\x[16][12] ), .ip2(n23656), .op(n23658) );
  or2_1 U27787 ( .ip1(n24079), .ip2(n23656), .op(n23657) );
  nand2_1 U27788 ( .ip1(n23658), .ip2(n23657), .op(n24437) );
  nor2_1 U27789 ( .ip1(n24371), .ip2(\x[16][11] ), .op(n23694) );
  inv_1 U27790 ( .ip(\x[16][9] ), .op(n23690) );
  inv_1 U27791 ( .ip(\x[16][8] ), .op(n23682) );
  nor2_1 U27792 ( .ip1(n23779), .ip2(n23682), .op(n23680) );
  inv_1 U27793 ( .ip(\x[16][6] ), .op(n23678) );
  nor2_1 U27794 ( .ip1(sig_in[6]), .ip2(n23678), .op(n23675) );
  inv_1 U27795 ( .ip(\x[16][4] ), .op(n23673) );
  and2_1 U27796 ( .ip1(n23659), .ip2(\x[16][2] ), .op(n23665) );
  nand2_1 U27797 ( .ip1(\x[16][1] ), .ip2(n20652), .op(n23663) );
  nand2_1 U27798 ( .ip1(\x[16][0] ), .ip2(n24143), .op(n23662) );
  nor2_1 U27799 ( .ip1(\x[16][2] ), .ip2(n23717), .op(n23661) );
  nor2_1 U27800 ( .ip1(\x[16][1] ), .ip2(n21685), .op(n23660) );
  not_ab_or_c_or_d U27801 ( .ip1(n23663), .ip2(n23662), .ip3(n23661), .ip4(
        n23660), .op(n23664) );
  not_ab_or_c_or_d U27802 ( .ip1(\x[16][3] ), .ip2(n24342), .ip3(n23665), 
        .ip4(n23664), .op(n23667) );
  nor2_1 U27803 ( .ip1(\x[16][3] ), .ip2(n24342), .op(n23666) );
  nor2_1 U27804 ( .ip1(n23667), .ip2(n23666), .op(n23668) );
  or2_1 U27805 ( .ip1(\x[16][4] ), .ip2(n23668), .op(n23670) );
  or2_1 U27806 ( .ip1(n23860), .ip2(n23668), .op(n23669) );
  nand2_1 U27807 ( .ip1(n23670), .ip2(n23669), .op(n23672) );
  nor2_1 U27808 ( .ip1(\x[16][5] ), .ip2(n24350), .op(n23671) );
  not_ab_or_c_or_d U27809 ( .ip1(sig_in[4]), .ip2(n23673), .ip3(n23672), .ip4(
        n23671), .op(n23674) );
  not_ab_or_c_or_d U27810 ( .ip1(\x[16][5] ), .ip2(n24482), .ip3(n23675), 
        .ip4(n23674), .op(n23677) );
  nor2_1 U27811 ( .ip1(\x[16][7] ), .ip2(n24044), .op(n23676) );
  not_ab_or_c_or_d U27812 ( .ip1(sig_in[6]), .ip2(n23678), .ip3(n23677), .ip4(
        n23676), .op(n23679) );
  not_ab_or_c_or_d U27813 ( .ip1(\x[16][7] ), .ip2(n24044), .ip3(n23680), 
        .ip4(n23679), .op(n23681) );
  or2_1 U27814 ( .ip1(sig_in[8]), .ip2(n23681), .op(n23684) );
  or2_1 U27815 ( .ip1(n23682), .ip2(n23681), .op(n23683) );
  nand2_1 U27816 ( .ip1(n23684), .ip2(n23683), .op(n23685) );
  or2_1 U27817 ( .ip1(\x[16][9] ), .ip2(n23685), .op(n23687) );
  or2_1 U27818 ( .ip1(n24043), .ip2(n23685), .op(n23686) );
  nand2_1 U27819 ( .ip1(n23687), .ip2(n23686), .op(n23689) );
  nor2_1 U27820 ( .ip1(\x[16][10] ), .ip2(n24370), .op(n23688) );
  not_ab_or_c_or_d U27821 ( .ip1(sig_in[9]), .ip2(n23690), .ip3(n23689), .ip4(
        n23688), .op(n23692) );
  and2_1 U27822 ( .ip1(n24370), .ip2(\x[16][10] ), .op(n23691) );
  not_ab_or_c_or_d U27823 ( .ip1(\x[16][11] ), .ip2(n24136), .ip3(n23692), 
        .ip4(n23691), .op(n23693) );
  nor2_1 U27824 ( .ip1(n23694), .ip2(n23693), .op(n24435) );
  inv_1 U27825 ( .ip(n24435), .op(n23695) );
  nand2_1 U27826 ( .ip1(n24437), .ip2(n23695), .op(n23700) );
  nor2_1 U27827 ( .ip1(\x[16][13] ), .ip2(n24137), .op(n23696) );
  or2_1 U27828 ( .ip1(sig_in[12]), .ip2(n23696), .op(n23699) );
  inv_1 U27829 ( .ip(\x[16][12] ), .op(n23697) );
  or2_1 U27830 ( .ip1(n23697), .ip2(n23696), .op(n23698) );
  nand2_1 U27831 ( .ip1(n23699), .ip2(n23698), .op(n24434) );
  nand2_1 U27832 ( .ip1(n23700), .ip2(n24434), .op(n23702) );
  nand2_1 U27833 ( .ip1(n24230), .ip2(\x[16][14] ), .op(n24436) );
  nor2_1 U27834 ( .ip1(\x[16][15] ), .ip2(n24090), .op(n24431) );
  inv_1 U27835 ( .ip(n24431), .op(n23705) );
  and2_1 U27836 ( .ip1(n24436), .ip2(n23705), .op(n23701) );
  nand2_1 U27837 ( .ip1(n23702), .ip2(n23701), .op(n23707) );
  or2_1 U27838 ( .ip1(n24382), .ip2(\x[16][14] ), .op(n23704) );
  nand2_1 U27839 ( .ip1(\x[16][15] ), .ip2(n24186), .op(n23703) );
  nand2_1 U27840 ( .ip1(n23704), .ip2(n23703), .op(n24433) );
  nand2_1 U27841 ( .ip1(n24433), .ip2(n23705), .op(n23706) );
  nand2_1 U27842 ( .ip1(n23707), .ip2(n23706), .op(n23708) );
  not_ab_or_c_or_d U27843 ( .ip1(n23711), .ip2(n23710), .ip3(n23709), .ip4(
        n23708), .op(n24722) );
  nor2_1 U27844 ( .ip1(n24384), .ip2(\x[18][15] ), .op(n23753) );
  inv_1 U27845 ( .ip(n23753), .op(n23801) );
  nand2_1 U27846 ( .ip1(\x[18][15] ), .ip2(n24186), .op(n24407) );
  or2_1 U27847 ( .ip1(n24382), .ip2(\x[18][14] ), .op(n23712) );
  nand2_1 U27848 ( .ip1(n24407), .ip2(n23712), .op(n24421) );
  nor2_1 U27849 ( .ip1(\x[17][15] ), .ip2(n24090), .op(n24429) );
  and2_1 U27850 ( .ip1(n24371), .ip2(\x[18][11] ), .op(n23747) );
  nor2_1 U27851 ( .ip1(\x[18][10] ), .ip2(n24457), .op(n23745) );
  nor2_1 U27852 ( .ip1(\x[18][9] ), .ip2(n24043), .op(n23739) );
  and2_1 U27853 ( .ip1(n23804), .ip2(\x[18][8] ), .op(n23737) );
  inv_1 U27854 ( .ip(\x[18][7] ), .op(n23734) );
  nor2_1 U27855 ( .ip1(n17732), .ip2(n23734), .op(n23731) );
  inv_1 U27856 ( .ip(\x[18][3] ), .op(n23720) );
  inv_1 U27857 ( .ip(\x[18][1] ), .op(n23714) );
  nor2_1 U27858 ( .ip1(sig_in[1]), .ip2(n23714), .op(n23716) );
  inv_1 U27859 ( .ip(\x[18][0] ), .op(n23713) );
  not_ab_or_c_or_d U27860 ( .ip1(n24467), .ip2(n23714), .ip3(sig_in[0]), .ip4(
        n23713), .op(n23715) );
  not_ab_or_c_or_d U27861 ( .ip1(\x[18][2] ), .ip2(n24470), .ip3(n23716), 
        .ip4(n23715), .op(n23719) );
  nor2_1 U27862 ( .ip1(\x[18][2] ), .ip2(n23717), .op(n23718) );
  not_ab_or_c_or_d U27863 ( .ip1(sig_in[3]), .ip2(n23720), .ip3(n23719), .ip4(
        n23718), .op(n23725) );
  nand2_1 U27864 ( .ip1(\x[18][5] ), .ip2(n24119), .op(n23723) );
  nand2_1 U27865 ( .ip1(\x[18][4] ), .ip2(n23721), .op(n23722) );
  nand2_1 U27866 ( .ip1(n23723), .ip2(n23722), .op(n23724) );
  not_ab_or_c_or_d U27867 ( .ip1(\x[18][3] ), .ip2(n22525), .ip3(n23725), 
        .ip4(n23724), .op(n23729) );
  nor2_1 U27868 ( .ip1(\x[18][6] ), .ip2(n24355), .op(n23728) );
  nor2_1 U27869 ( .ip1(\x[18][5] ), .ip2(n24350), .op(n23727) );
  not_ab_or_c_or_d U27870 ( .ip1(\x[18][5] ), .ip2(n24482), .ip3(\x[18][4] ), 
        .ip4(n24256), .op(n23726) );
  nor4_1 U27871 ( .ip1(n23729), .ip2(n23728), .ip3(n23727), .ip4(n23726), .op(
        n23730) );
  not_ab_or_c_or_d U27872 ( .ip1(\x[18][6] ), .ip2(n24355), .ip3(n23731), 
        .ip4(n23730), .op(n23733) );
  nor2_1 U27873 ( .ip1(\x[18][8] ), .ip2(n23971), .op(n23732) );
  not_ab_or_c_or_d U27874 ( .ip1(sig_in[7]), .ip2(n23734), .ip3(n23733), .ip4(
        n23732), .op(n23736) );
  and2_1 U27875 ( .ip1(n24043), .ip2(\x[18][9] ), .op(n23735) );
  nor3_1 U27876 ( .ip1(n23737), .ip2(n23736), .ip3(n23735), .op(n23738) );
  nor2_1 U27877 ( .ip1(n23739), .ip2(n23738), .op(n23740) );
  or2_1 U27878 ( .ip1(\x[18][10] ), .ip2(n23740), .op(n23742) );
  or2_1 U27879 ( .ip1(n24457), .ip2(n23740), .op(n23741) );
  nand2_1 U27880 ( .ip1(n23742), .ip2(n23741), .op(n23744) );
  nor2_1 U27881 ( .ip1(\x[18][11] ), .ip2(n24239), .op(n23743) );
  nor3_1 U27882 ( .ip1(n23745), .ip2(n23744), .ip3(n23743), .op(n23746) );
  nor2_1 U27883 ( .ip1(n23747), .ip2(n23746), .op(n24422) );
  nand2_1 U27884 ( .ip1(\x[18][12] ), .ip2(n24233), .op(n24405) );
  nand2_1 U27885 ( .ip1(n24422), .ip2(n24405), .op(n23752) );
  nor2_1 U27886 ( .ip1(\x[18][13] ), .ip2(n24137), .op(n23748) );
  or2_1 U27887 ( .ip1(sig_in[12]), .ip2(n23748), .op(n23751) );
  inv_1 U27888 ( .ip(\x[18][12] ), .op(n23749) );
  or2_1 U27889 ( .ip1(n23749), .ip2(n23748), .op(n23750) );
  nand2_1 U27890 ( .ip1(n23751), .ip2(n23750), .op(n24419) );
  nand2_1 U27891 ( .ip1(n23752), .ip2(n24419), .op(n23755) );
  and2_1 U27892 ( .ip1(n24332), .ip2(\x[18][13] ), .op(n23754) );
  not_ab_or_c_or_d U27893 ( .ip1(\x[18][14] ), .ip2(n23938), .ip3(n23754), 
        .ip4(n23753), .op(n24406) );
  nand2_1 U27894 ( .ip1(n23755), .ip2(n24406), .op(n23799) );
  and2_1 U27895 ( .ip1(n24461), .ip2(\x[17][7] ), .op(n23769) );
  inv_1 U27896 ( .ip(\x[17][4] ), .op(n23767) );
  nor2_1 U27897 ( .ip1(n24462), .ip2(n23767), .op(n23764) );
  inv_1 U27898 ( .ip(n24342), .op(n24251) );
  inv_1 U27899 ( .ip(\x[17][3] ), .op(n23762) );
  nor2_1 U27900 ( .ip1(\x[17][2] ), .ip2(n24463), .op(n23761) );
  inv_1 U27901 ( .ip(\x[17][1] ), .op(n23757) );
  nor2_1 U27902 ( .ip1(n24464), .ip2(n23757), .op(n23759) );
  inv_1 U27903 ( .ip(\x[17][0] ), .op(n23756) );
  not_ab_or_c_or_d U27904 ( .ip1(n24467), .ip2(n23757), .ip3(sig_in[0]), .ip4(
        n23756), .op(n23758) );
  not_ab_or_c_or_d U27905 ( .ip1(\x[17][2] ), .ip2(n24470), .ip3(n23759), 
        .ip4(n23758), .op(n23760) );
  not_ab_or_c_or_d U27906 ( .ip1(n24251), .ip2(n23762), .ip3(n23761), .ip4(
        n23760), .op(n23763) );
  not_ab_or_c_or_d U27907 ( .ip1(\x[17][3] ), .ip2(n24342), .ip3(n23764), 
        .ip4(n23763), .op(n23766) );
  nor2_1 U27908 ( .ip1(\x[17][5] ), .ip2(n24350), .op(n23765) );
  not_ab_or_c_or_d U27909 ( .ip1(sig_in[4]), .ip2(n23767), .ip3(n23766), .ip4(
        n23765), .op(n23768) );
  not_ab_or_c_or_d U27910 ( .ip1(\x[17][5] ), .ip2(n24482), .ip3(n23769), 
        .ip4(n23768), .op(n23774) );
  nand2_1 U27911 ( .ip1(\x[17][6] ), .ip2(n24485), .op(n23773) );
  nor2_1 U27912 ( .ip1(\x[17][7] ), .ip2(n24044), .op(n23772) );
  not_ab_or_c_or_d U27913 ( .ip1(\x[17][7] ), .ip2(n24044), .ip3(\x[17][6] ), 
        .ip4(n23770), .op(n23771) );
  not_ab_or_c_or_d U27914 ( .ip1(n23774), .ip2(n23773), .ip3(n23772), .ip4(
        n23771), .op(n23775) );
  nand2_1 U27915 ( .ip1(\x[17][8] ), .ip2(n23775), .op(n23778) );
  nor2_1 U27916 ( .ip1(\x[17][9] ), .ip2(n24164), .op(n23777) );
  nor2_1 U27917 ( .ip1(\x[17][8] ), .ip2(n23775), .op(n23776) );
  ab_or_c_or_d U27918 ( .ip1(n23779), .ip2(n23778), .ip3(n23777), .ip4(n23776), 
        .op(n23783) );
  nand2_1 U27919 ( .ip1(\x[17][10] ), .ip2(n24370), .op(n23782) );
  nand2_1 U27920 ( .ip1(\x[17][11] ), .ip2(n24239), .op(n23781) );
  nand2_1 U27921 ( .ip1(\x[17][9] ), .ip2(n24269), .op(n23780) );
  and4_1 U27922 ( .ip1(n23783), .ip2(n23782), .ip3(n23781), .ip4(n23780), .op(
        n23787) );
  nor2_1 U27923 ( .ip1(n24239), .ip2(\x[17][11] ), .op(n23785) );
  not_ab_or_c_or_d U27924 ( .ip1(\x[17][11] ), .ip2(n24136), .ip3(\x[17][10] ), 
        .ip4(n23980), .op(n23784) );
  or2_1 U27925 ( .ip1(n23785), .ip2(n23784), .op(n23786) );
  nor2_1 U27926 ( .ip1(n23787), .ip2(n23786), .op(n24441) );
  nor2_1 U27927 ( .ip1(\x[17][13] ), .ip2(n24376), .op(n23788) );
  or2_1 U27928 ( .ip1(sig_in[12]), .ip2(n23788), .op(n23791) );
  inv_1 U27929 ( .ip(\x[17][12] ), .op(n23789) );
  or2_1 U27930 ( .ip1(n23789), .ip2(n23788), .op(n23790) );
  nand2_1 U27931 ( .ip1(n23791), .ip2(n23790), .op(n24428) );
  or2_1 U27932 ( .ip1(n24382), .ip2(\x[17][14] ), .op(n23792) );
  nand3_1 U27933 ( .ip1(n24441), .ip2(n24428), .ip3(n23792), .op(n23796) );
  and2_1 U27934 ( .ip1(n24235), .ip2(\x[17][13] ), .op(n23793) );
  or2_1 U27935 ( .ip1(\x[17][12] ), .ip2(n23793), .op(n23795) );
  or2_1 U27936 ( .ip1(n24079), .ip2(n23793), .op(n23794) );
  nand2_1 U27937 ( .ip1(n23795), .ip2(n23794), .op(n24444) );
  nand2_1 U27938 ( .ip1(\x[17][14] ), .ip2(n23938), .op(n24426) );
  nand3_1 U27939 ( .ip1(n23796), .ip2(n24444), .ip3(n24426), .op(n23797) );
  nand2_1 U27940 ( .ip1(\x[17][15] ), .ip2(n24186), .op(n24446) );
  nand2_1 U27941 ( .ip1(n23797), .ip2(n24446), .op(n23798) );
  nand2_1 U27942 ( .ip1(n23799), .ip2(n23798), .op(n23800) );
  not_ab_or_c_or_d U27943 ( .ip1(n23801), .ip2(n24421), .ip3(n24429), .ip4(
        n23800), .op(n24701) );
  and2_1 U27944 ( .ip1(n24081), .ip2(\x[19][13] ), .op(n23802) );
  nor2_1 U27945 ( .ip1(\x[19][15] ), .ip2(n24090), .op(n24414) );
  not_ab_or_c_or_d U27946 ( .ip1(\x[19][14] ), .ip2(n23938), .ip3(n23802), 
        .ip4(n24414), .op(n24410) );
  nand2_1 U27947 ( .ip1(\x[19][12] ), .ip2(n24449), .op(n23803) );
  nand2_1 U27948 ( .ip1(n24410), .ip2(n23803), .op(n24409) );
  nand2_1 U27949 ( .ip1(\x[19][15] ), .ip2(n24186), .op(n23894) );
  inv_1 U27950 ( .ip(\x[19][11] ), .op(n23834) );
  and2_1 U27951 ( .ip1(n24451), .ip2(\x[19][10] ), .op(n23831) );
  inv_1 U27952 ( .ip(\x[19][9] ), .op(n23829) );
  and2_1 U27953 ( .ip1(n23804), .ip2(\x[19][8] ), .op(n23826) );
  inv_1 U27954 ( .ip(\x[19][6] ), .op(n23824) );
  nor2_1 U27955 ( .ip1(\x[19][5] ), .ip2(n24350), .op(n23818) );
  and2_1 U27956 ( .ip1(n23721), .ip2(\x[19][4] ), .op(n23816) );
  inv_1 U27957 ( .ip(\x[19][3] ), .op(n23813) );
  and2_1 U27958 ( .ip1(n24335), .ip2(\x[19][2] ), .op(n23810) );
  nand2_1 U27959 ( .ip1(\x[19][1] ), .ip2(n20652), .op(n23808) );
  nand2_1 U27960 ( .ip1(\x[19][0] ), .ip2(n24143), .op(n23807) );
  nor2_1 U27961 ( .ip1(\x[19][2] ), .ip2(n24463), .op(n23806) );
  nor2_1 U27962 ( .ip1(\x[19][1] ), .ip2(n20652), .op(n23805) );
  not_ab_or_c_or_d U27963 ( .ip1(n23808), .ip2(n23807), .ip3(n23806), .ip4(
        n23805), .op(n23809) );
  not_ab_or_c_or_d U27964 ( .ip1(\x[19][3] ), .ip2(n24342), .ip3(n23810), 
        .ip4(n23809), .op(n23812) );
  nor2_1 U27965 ( .ip1(\x[19][4] ), .ip2(n24347), .op(n23811) );
  not_ab_or_c_or_d U27966 ( .ip1(n23251), .ip2(n23813), .ip3(n23812), .ip4(
        n23811), .op(n23815) );
  and2_1 U27967 ( .ip1(n24350), .ip2(\x[19][5] ), .op(n23814) );
  nor3_1 U27968 ( .ip1(n23816), .ip2(n23815), .ip3(n23814), .op(n23817) );
  nor2_1 U27969 ( .ip1(n23818), .ip2(n23817), .op(n23819) );
  or2_1 U27970 ( .ip1(\x[19][6] ), .ip2(n23819), .op(n23821) );
  or2_1 U27971 ( .ip1(n23770), .ip2(n23819), .op(n23820) );
  nand2_1 U27972 ( .ip1(n23821), .ip2(n23820), .op(n23823) );
  nor2_1 U27973 ( .ip1(\x[19][7] ), .ip2(n24492), .op(n23822) );
  not_ab_or_c_or_d U27974 ( .ip1(sig_in[6]), .ip2(n23824), .ip3(n23823), .ip4(
        n23822), .op(n23825) );
  not_ab_or_c_or_d U27975 ( .ip1(\x[19][7] ), .ip2(n24142), .ip3(n23826), 
        .ip4(n23825), .op(n23828) );
  nor2_1 U27976 ( .ip1(\x[19][8] ), .ip2(n23971), .op(n23827) );
  not_ab_or_c_or_d U27977 ( .ip1(sig_in[9]), .ip2(n23829), .ip3(n23828), .ip4(
        n23827), .op(n23830) );
  not_ab_or_c_or_d U27978 ( .ip1(\x[19][9] ), .ip2(n24269), .ip3(n23831), 
        .ip4(n23830), .op(n23833) );
  nor2_1 U27979 ( .ip1(\x[19][10] ), .ip2(n24457), .op(n23832) );
  not_ab_or_c_or_d U27980 ( .ip1(sig_in[11]), .ip2(n23834), .ip3(n23833), 
        .ip4(n23832), .op(n23835) );
  or2_1 U27981 ( .ip1(\x[19][11] ), .ip2(n23835), .op(n23837) );
  or2_1 U27982 ( .ip1(n24136), .ip2(n23835), .op(n23836) );
  nand2_1 U27983 ( .ip1(n23837), .ip2(n23836), .op(n24418) );
  nor2_1 U27984 ( .ip1(\x[19][13] ), .ip2(n24081), .op(n23839) );
  nor2_1 U27985 ( .ip1(\x[19][12] ), .ip2(n24450), .op(n23838) );
  or2_1 U27986 ( .ip1(n23839), .ip2(n23838), .op(n24411) );
  or2_1 U27987 ( .ip1(n24185), .ip2(\x[19][14] ), .op(n23840) );
  nand2_1 U27988 ( .ip1(n23894), .ip2(n23840), .op(n24412) );
  nor3_1 U27989 ( .ip1(n24418), .ip2(n24411), .ip3(n24412), .op(n23893) );
  and2_1 U27990 ( .ip1(n24235), .ip2(\x[20][13] ), .op(n23841) );
  or2_1 U27991 ( .ip1(\x[20][12] ), .ip2(n23841), .op(n23843) );
  or2_1 U27992 ( .ip1(n24449), .ip2(n23841), .op(n23842) );
  nand2_1 U27993 ( .ip1(n23843), .ip2(n23842), .op(n24389) );
  and2_1 U27994 ( .ip1(n24461), .ip2(\x[20][7] ), .op(n23865) );
  inv_1 U27995 ( .ip(\x[20][5] ), .op(n23863) );
  nor2_1 U27996 ( .ip1(sig_in[5]), .ip2(n23863), .op(n23859) );
  inv_1 U27997 ( .ip(\x[20][3] ), .op(n23850) );
  inv_1 U27998 ( .ip(\x[20][1] ), .op(n23845) );
  nor2_1 U27999 ( .ip1(sig_in[1]), .ip2(n23845), .op(n23847) );
  inv_1 U28000 ( .ip(\x[20][0] ), .op(n23844) );
  not_ab_or_c_or_d U28001 ( .ip1(n24467), .ip2(n23845), .ip3(sig_in[0]), .ip4(
        n23844), .op(n23846) );
  not_ab_or_c_or_d U28002 ( .ip1(\x[20][2] ), .ip2(n24470), .ip3(n23847), 
        .ip4(n23846), .op(n23849) );
  nor2_1 U28003 ( .ip1(\x[20][2] ), .ip2(n24463), .op(n23848) );
  not_ab_or_c_or_d U28004 ( .ip1(n24251), .ip2(n23850), .ip3(n23849), .ip4(
        n23848), .op(n23851) );
  or2_1 U28005 ( .ip1(\x[20][3] ), .ip2(n23851), .op(n23853) );
  or2_1 U28006 ( .ip1(n22795), .ip2(n23851), .op(n23852) );
  nand2_1 U28007 ( .ip1(n23853), .ip2(n23852), .op(n23854) );
  or2_1 U28008 ( .ip1(sig_in[4]), .ip2(n23854), .op(n23857) );
  inv_1 U28009 ( .ip(\x[20][4] ), .op(n23855) );
  or2_1 U28010 ( .ip1(n23855), .ip2(n23854), .op(n23856) );
  nand2_1 U28011 ( .ip1(n23857), .ip2(n23856), .op(n23858) );
  not_ab_or_c_or_d U28012 ( .ip1(\x[20][4] ), .ip2(n23860), .ip3(n23859), 
        .ip4(n23858), .op(n23862) );
  nor2_1 U28013 ( .ip1(\x[20][6] ), .ip2(n24355), .op(n23861) );
  not_ab_or_c_or_d U28014 ( .ip1(sig_in[5]), .ip2(n23863), .ip3(n23862), .ip4(
        n23861), .op(n23864) );
  not_ab_or_c_or_d U28015 ( .ip1(\x[20][6] ), .ip2(n24045), .ip3(n23865), 
        .ip4(n23864), .op(n23868) );
  nor2_1 U28016 ( .ip1(\x[20][9] ), .ip2(n24269), .op(n23869) );
  nor2_1 U28017 ( .ip1(\x[20][8] ), .ip2(n23971), .op(n23867) );
  nor2_1 U28018 ( .ip1(\x[20][7] ), .ip2(n24492), .op(n23866) );
  nor4_1 U28019 ( .ip1(n23868), .ip2(n23869), .ip3(n23867), .ip4(n23866), .op(
        n23875) );
  nand2_1 U28020 ( .ip1(n24370), .ip2(\x[20][10] ), .op(n23873) );
  inv_1 U28021 ( .ip(n23869), .op(n23870) );
  nand3_1 U28022 ( .ip1(\x[20][8] ), .ip2(n23971), .ip3(n23870), .op(n23872)
         );
  nand2_1 U28023 ( .ip1(\x[20][11] ), .ip2(n24371), .op(n23871) );
  nand3_1 U28024 ( .ip1(n23873), .ip2(n23872), .ip3(n23871), .op(n23874) );
  not_ab_or_c_or_d U28025 ( .ip1(\x[20][9] ), .ip2(n24455), .ip3(n23875), 
        .ip4(n23874), .op(n23879) );
  nor2_1 U28026 ( .ip1(n21793), .ip2(\x[20][11] ), .op(n23877) );
  not_ab_or_c_or_d U28027 ( .ip1(\x[20][11] ), .ip2(n24136), .ip3(\x[20][10] ), 
        .ip4(n24370), .op(n23876) );
  or2_1 U28028 ( .ip1(n23877), .ip2(n23876), .op(n23878) );
  nor2_1 U28029 ( .ip1(n23879), .ip2(n23878), .op(n24401) );
  inv_1 U28030 ( .ip(n24401), .op(n23880) );
  nand2_1 U28031 ( .ip1(n24389), .ip2(n23880), .op(n23885) );
  nor2_1 U28032 ( .ip1(\x[20][13] ), .ip2(n24081), .op(n23881) );
  or2_1 U28033 ( .ip1(sig_in[12]), .ip2(n23881), .op(n23884) );
  inv_1 U28034 ( .ip(\x[20][12] ), .op(n23882) );
  or2_1 U28035 ( .ip1(n23882), .ip2(n23881), .op(n23883) );
  nand2_1 U28036 ( .ip1(n23884), .ip2(n23883), .op(n24400) );
  nand2_1 U28037 ( .ip1(n23885), .ip2(n24400), .op(n23887) );
  nor2_1 U28038 ( .ip1(\x[20][15] ), .ip2(n24090), .op(n24395) );
  inv_1 U28039 ( .ip(n24395), .op(n23889) );
  nand2_1 U28040 ( .ip1(n23938), .ip2(\x[20][14] ), .op(n24388) );
  and2_1 U28041 ( .ip1(n23889), .ip2(n24388), .op(n23886) );
  nand2_1 U28042 ( .ip1(n23887), .ip2(n23886), .op(n23891) );
  nand2_1 U28043 ( .ip1(\x[20][15] ), .ip2(n24186), .op(n24390) );
  or2_1 U28044 ( .ip1(n24382), .ip2(\x[20][14] ), .op(n23888) );
  nand2_1 U28045 ( .ip1(n24390), .ip2(n23888), .op(n24398) );
  nand2_1 U28046 ( .ip1(n23889), .ip2(n24398), .op(n23890) );
  nand2_1 U28047 ( .ip1(n23891), .ip2(n23890), .op(n23892) );
  not_ab_or_c_or_d U28048 ( .ip1(n24409), .ip2(n23894), .ip3(n23893), .ip4(
        n23892), .op(n24790) );
  and2_1 U28049 ( .ip1(n23895), .ip2(\x[23][13] ), .op(n23896) );
  nor2_1 U28050 ( .ip1(\x[23][15] ), .ip2(n24090), .op(n23903) );
  not_ab_or_c_or_d U28051 ( .ip1(\x[23][14] ), .ip2(n24327), .ip3(n23896), 
        .ip4(n23903), .op(n23996) );
  nor2_1 U28052 ( .ip1(\x[23][13] ), .ip2(n24081), .op(n23898) );
  nor2_1 U28053 ( .ip1(\x[23][12] ), .ip2(n24079), .op(n23897) );
  nor2_1 U28054 ( .ip1(n23898), .ip2(n23897), .op(n24315) );
  inv_1 U28055 ( .ip(n24315), .op(n23995) );
  nand2_1 U28056 ( .ip1(n24329), .ip2(\x[23][15] ), .op(n24308) );
  inv_1 U28057 ( .ip(n24308), .op(n23899) );
  or2_1 U28058 ( .ip1(sig_in[14]), .ip2(n23899), .op(n23902) );
  inv_1 U28059 ( .ip(\x[23][14] ), .op(n23900) );
  or2_1 U28060 ( .ip1(n23900), .ip2(n23899), .op(n23901) );
  nand2_1 U28061 ( .ip1(n23902), .ip2(n23901), .op(n24314) );
  nor2_1 U28062 ( .ip1(n23903), .ip2(n24314), .op(n23994) );
  nor2_1 U28063 ( .ip1(n24456), .ip2(\x[23][11] ), .op(n23935) );
  nor2_1 U28064 ( .ip1(\x[23][9] ), .ip2(n24164), .op(n23925) );
  inv_1 U28065 ( .ip(\x[23][8] ), .op(n23904) );
  nor3_1 U28066 ( .ip1(n23779), .ip2(n23925), .ip3(n23904), .op(n23927) );
  nor2_1 U28067 ( .ip1(\x[23][8] ), .ip2(n24100), .op(n23924) );
  nor2_1 U28068 ( .ip1(\x[23][7] ), .ip2(n24492), .op(n23923) );
  and2_1 U28069 ( .ip1(n24461), .ip2(\x[23][7] ), .op(n23919) );
  nor3_1 U28070 ( .ip1(n24045), .ip2(\x[23][6] ), .ip3(n23919), .op(n23921) );
  nor2_1 U28071 ( .ip1(\x[23][5] ), .ip2(n24350), .op(n23914) );
  inv_1 U28072 ( .ip(\x[23][4] ), .op(n23905) );
  nor3_1 U28073 ( .ip1(n24462), .ip2(n23914), .ip3(n23905), .op(n23917) );
  and2_1 U28074 ( .ip1(n24335), .ip2(\x[23][2] ), .op(n23911) );
  nand2_1 U28075 ( .ip1(\x[23][1] ), .ip2(n21685), .op(n23909) );
  nand2_1 U28076 ( .ip1(\x[23][0] ), .ip2(n24143), .op(n23908) );
  nor2_1 U28077 ( .ip1(\x[23][2] ), .ip2(n24463), .op(n23907) );
  nor2_1 U28078 ( .ip1(\x[23][1] ), .ip2(n21685), .op(n23906) );
  not_ab_or_c_or_d U28079 ( .ip1(n23909), .ip2(n23908), .ip3(n23907), .ip4(
        n23906), .op(n23910) );
  not_ab_or_c_or_d U28080 ( .ip1(\x[23][3] ), .ip2(n24342), .ip3(n23911), 
        .ip4(n23910), .op(n23915) );
  nor2_1 U28081 ( .ip1(\x[23][3] ), .ip2(n24342), .op(n23913) );
  nor2_1 U28082 ( .ip1(\x[23][4] ), .ip2(n23860), .op(n23912) );
  nor4_1 U28083 ( .ip1(n23915), .ip2(n23914), .ip3(n23913), .ip4(n23912), .op(
        n23916) );
  ab_or_c_or_d U28084 ( .ip1(\x[23][5] ), .ip2(n24119), .ip3(n23917), .ip4(
        n23916), .op(n23918) );
  not_ab_or_c_or_d U28085 ( .ip1(\x[23][6] ), .ip2(n24485), .ip3(n23919), 
        .ip4(n23918), .op(n23920) );
  or2_1 U28086 ( .ip1(n23921), .ip2(n23920), .op(n23922) );
  nor4_1 U28087 ( .ip1(n23925), .ip2(n23924), .ip3(n23923), .ip4(n23922), .op(
        n23926) );
  not_ab_or_c_or_d U28088 ( .ip1(\x[23][9] ), .ip2(n24269), .ip3(n23927), 
        .ip4(n23926), .op(n23928) );
  or2_1 U28089 ( .ip1(sig_in[10]), .ip2(n23928), .op(n23930) );
  inv_1 U28090 ( .ip(\x[23][10] ), .op(n23931) );
  or2_1 U28091 ( .ip1(n23931), .ip2(n23928), .op(n23929) );
  nand2_1 U28092 ( .ip1(n23930), .ip2(n23929), .op(n23933) );
  nor2_1 U28093 ( .ip1(sig_in[10]), .ip2(n23931), .op(n23932) );
  not_ab_or_c_or_d U28094 ( .ip1(\x[23][11] ), .ip2(n24136), .ip3(n23933), 
        .ip4(n23932), .op(n23934) );
  nor2_1 U28095 ( .ip1(n23935), .ip2(n23934), .op(n24316) );
  nand2_1 U28096 ( .ip1(\x[23][12] ), .ip2(n24233), .op(n23936) );
  nand2_1 U28097 ( .ip1(n23996), .ip2(n23936), .op(n24309) );
  or2_1 U28098 ( .ip1(n24316), .ip2(n24309), .op(n23992) );
  and2_1 U28099 ( .ip1(n24081), .ip2(\x[22][13] ), .op(n23937) );
  nor2_1 U28100 ( .ip1(\x[22][15] ), .ip2(n24090), .op(n23942) );
  not_ab_or_c_or_d U28101 ( .ip1(\x[22][14] ), .ip2(n24327), .ip3(n23937), 
        .ip4(n23942), .op(n24325) );
  nand2_1 U28102 ( .ip1(\x[22][12] ), .ip2(n24450), .op(n24322) );
  nand2_1 U28103 ( .ip1(n24325), .ip2(n24322), .op(n23943) );
  nor2_1 U28104 ( .ip1(\x[22][14] ), .ip2(n23938), .op(n23939) );
  or2_1 U28105 ( .ip1(\x[22][15] ), .ip2(n23939), .op(n23941) );
  or2_1 U28106 ( .ip1(n24329), .ip2(n23939), .op(n23940) );
  nand2_1 U28107 ( .ip1(n23941), .ip2(n23940), .op(n23989) );
  or2_1 U28108 ( .ip1(n23942), .ip2(n23989), .op(n24386) );
  nand2_1 U28109 ( .ip1(n23943), .ip2(n24386), .op(n23991) );
  nor2_1 U28110 ( .ip1(\x[22][13] ), .ip2(n24137), .op(n23944) );
  or2_1 U28111 ( .ip1(sig_in[12]), .ip2(n23944), .op(n23947) );
  inv_1 U28112 ( .ip(\x[22][12] ), .op(n23945) );
  or2_1 U28113 ( .ip1(n23945), .ip2(n23944), .op(n23946) );
  nand2_1 U28114 ( .ip1(n23947), .ip2(n23946), .op(n24323) );
  nor2_1 U28115 ( .ip1(\x[22][10] ), .ip2(n24457), .op(n23948) );
  or2_1 U28116 ( .ip1(sig_in[11]), .ip2(n23948), .op(n23951) );
  inv_1 U28117 ( .ip(\x[22][11] ), .op(n23949) );
  or2_1 U28118 ( .ip1(n23949), .ip2(n23948), .op(n23950) );
  nand2_1 U28119 ( .ip1(n23951), .ip2(n23950), .op(n23986) );
  inv_1 U28120 ( .ip(\x[22][7] ), .op(n23974) );
  nor2_1 U28121 ( .ip1(n17732), .ip2(n23974), .op(n23970) );
  inv_1 U28122 ( .ip(\x[22][5] ), .op(n23968) );
  nor2_1 U28123 ( .ip1(sig_in[5]), .ip2(n23968), .op(n23965) );
  inv_1 U28124 ( .ip(\x[22][3] ), .op(n23963) );
  and2_1 U28125 ( .ip1(n24107), .ip2(\x[22][2] ), .op(n23960) );
  inv_1 U28126 ( .ip(\x[22][1] ), .op(n23953) );
  inv_1 U28127 ( .ip(\x[22][0] ), .op(n23952) );
  not_ab_or_c_or_d U28128 ( .ip1(n24467), .ip2(n23953), .ip3(sig_in[0]), .ip4(
        n23952), .op(n23954) );
  or2_1 U28129 ( .ip1(\x[22][1] ), .ip2(n23954), .op(n23956) );
  or2_1 U28130 ( .ip1(n20652), .ip2(n23954), .op(n23955) );
  nand2_1 U28131 ( .ip1(n23956), .ip2(n23955), .op(n23958) );
  nor2_1 U28132 ( .ip1(\x[22][2] ), .ip2(n24463), .op(n23957) );
  nor2_1 U28133 ( .ip1(n23958), .ip2(n23957), .op(n23959) );
  not_ab_or_c_or_d U28134 ( .ip1(\x[22][3] ), .ip2(n22795), .ip3(n23960), 
        .ip4(n23959), .op(n23962) );
  nor2_1 U28135 ( .ip1(\x[22][4] ), .ip2(n24347), .op(n23961) );
  not_ab_or_c_or_d U28136 ( .ip1(n24251), .ip2(n23963), .ip3(n23962), .ip4(
        n23961), .op(n23964) );
  not_ab_or_c_or_d U28137 ( .ip1(\x[22][4] ), .ip2(n24256), .ip3(n23965), 
        .ip4(n23964), .op(n23967) );
  nor2_1 U28138 ( .ip1(\x[22][6] ), .ip2(n24355), .op(n23966) );
  not_ab_or_c_or_d U28139 ( .ip1(sig_in[5]), .ip2(n23968), .ip3(n23967), .ip4(
        n23966), .op(n23969) );
  not_ab_or_c_or_d U28140 ( .ip1(\x[22][6] ), .ip2(n24045), .ip3(n23970), 
        .ip4(n23969), .op(n23973) );
  nor2_1 U28141 ( .ip1(\x[22][8] ), .ip2(n23971), .op(n23972) );
  not_ab_or_c_or_d U28142 ( .ip1(sig_in[7]), .ip2(n23974), .ip3(n23973), .ip4(
        n23972), .op(n23975) );
  or2_1 U28143 ( .ip1(\x[22][8] ), .ip2(n23975), .op(n23977) );
  or2_1 U28144 ( .ip1(n24491), .ip2(n23975), .op(n23976) );
  nand2_1 U28145 ( .ip1(n23977), .ip2(n23976), .op(n23979) );
  nor2_1 U28146 ( .ip1(\x[22][9] ), .ip2(n24164), .op(n23978) );
  or2_1 U28147 ( .ip1(n23979), .ip2(n23978), .op(n23984) );
  nand2_1 U28148 ( .ip1(\x[22][10] ), .ip2(n23980), .op(n23983) );
  nand2_1 U28149 ( .ip1(\x[22][9] ), .ip2(n23981), .op(n23982) );
  nand3_1 U28150 ( .ip1(n23984), .ip2(n23983), .ip3(n23982), .op(n23985) );
  nand2_1 U28151 ( .ip1(n23986), .ip2(n23985), .op(n23988) );
  nand2_1 U28152 ( .ip1(\x[22][11] ), .ip2(n24239), .op(n23987) );
  nand2_1 U28153 ( .ip1(n23988), .ip2(n23987), .op(n24320) );
  nand3_1 U28154 ( .ip1(n23989), .ip2(n24323), .ip3(n24320), .op(n23990) );
  nand3_1 U28155 ( .ip1(n23992), .ip2(n23991), .ip3(n23990), .op(n23993) );
  not_ab_or_c_or_d U28156 ( .ip1(n23996), .ip2(n23995), .ip3(n23994), .ip4(
        n23993), .op(n24793) );
  nor2_1 U28157 ( .ip1(\x[24][14] ), .ip2(n24327), .op(n23997) );
  or2_1 U28158 ( .ip1(\x[24][15] ), .ip2(n23997), .op(n23999) );
  or2_1 U28159 ( .ip1(n23143), .ip2(n23997), .op(n23998) );
  nand2_1 U28160 ( .ip1(n23999), .ip2(n23998), .op(n24301) );
  nor2_1 U28161 ( .ip1(\x[24][13] ), .ip2(n24137), .op(n24000) );
  or2_1 U28162 ( .ip1(sig_in[12]), .ip2(n24000), .op(n24003) );
  inv_1 U28163 ( .ip(\x[24][12] ), .op(n24001) );
  or2_1 U28164 ( .ip1(n24001), .ip2(n24000), .op(n24002) );
  nand2_1 U28165 ( .ip1(n24003), .ip2(n24002), .op(n24305) );
  inv_1 U28166 ( .ip(\x[24][11] ), .op(n24035) );
  nor2_1 U28167 ( .ip1(n24035), .ip2(n17981), .op(n24037) );
  and2_1 U28168 ( .ip1(n24451), .ip2(\x[24][10] ), .op(n24032) );
  inv_1 U28169 ( .ip(\x[24][9] ), .op(n24030) );
  nor2_1 U28170 ( .ip1(\x[24][8] ), .ip2(n24100), .op(n24029) );
  inv_1 U28171 ( .ip(\x[24][7] ), .op(n24022) );
  nor2_1 U28172 ( .ip1(n17732), .ip2(n24022), .op(n24020) );
  inv_1 U28173 ( .ip(\x[24][3] ), .op(n24010) );
  inv_1 U28174 ( .ip(\x[24][1] ), .op(n24005) );
  nor2_1 U28175 ( .ip1(n24464), .ip2(n24005), .op(n24007) );
  inv_1 U28176 ( .ip(\x[24][0] ), .op(n24004) );
  not_ab_or_c_or_d U28177 ( .ip1(n24467), .ip2(n24005), .ip3(sig_in[0]), .ip4(
        n24004), .op(n24006) );
  not_ab_or_c_or_d U28178 ( .ip1(\x[24][2] ), .ip2(n24470), .ip3(n24007), 
        .ip4(n24006), .op(n24009) );
  nor2_1 U28179 ( .ip1(\x[24][2] ), .ip2(n24463), .op(n24008) );
  not_ab_or_c_or_d U28180 ( .ip1(n24251), .ip2(n24010), .ip3(n24009), .ip4(
        n24008), .op(n24014) );
  nand2_1 U28181 ( .ip1(\x[24][5] ), .ip2(n24119), .op(n24012) );
  nand2_1 U28182 ( .ip1(\x[24][4] ), .ip2(n23860), .op(n24011) );
  nand2_1 U28183 ( .ip1(n24012), .ip2(n24011), .op(n24013) );
  not_ab_or_c_or_d U28184 ( .ip1(\x[24][3] ), .ip2(n22795), .ip3(n24014), 
        .ip4(n24013), .op(n24018) );
  nor2_1 U28185 ( .ip1(\x[24][5] ), .ip2(n24350), .op(n24017) );
  nor2_1 U28186 ( .ip1(\x[24][6] ), .ip2(n24355), .op(n24016) );
  not_ab_or_c_or_d U28187 ( .ip1(\x[24][5] ), .ip2(n24482), .ip3(\x[24][4] ), 
        .ip4(n24256), .op(n24015) );
  nor4_1 U28188 ( .ip1(n24018), .ip2(n24017), .ip3(n24016), .ip4(n24015), .op(
        n24019) );
  not_ab_or_c_or_d U28189 ( .ip1(\x[24][6] ), .ip2(n24045), .ip3(n24020), 
        .ip4(n24019), .op(n24021) );
  or2_1 U28190 ( .ip1(sig_in[7]), .ip2(n24021), .op(n24024) );
  or2_1 U28191 ( .ip1(n24022), .ip2(n24021), .op(n24023) );
  nand2_1 U28192 ( .ip1(n24024), .ip2(n24023), .op(n24025) );
  or2_1 U28193 ( .ip1(\x[24][8] ), .ip2(n24025), .op(n24027) );
  or2_1 U28194 ( .ip1(n24491), .ip2(n24025), .op(n24026) );
  nand2_1 U28195 ( .ip1(n24027), .ip2(n24026), .op(n24028) );
  not_ab_or_c_or_d U28196 ( .ip1(sig_in[9]), .ip2(n24030), .ip3(n24029), .ip4(
        n24028), .op(n24031) );
  not_ab_or_c_or_d U28197 ( .ip1(\x[24][9] ), .ip2(n24269), .ip3(n24032), 
        .ip4(n24031), .op(n24034) );
  nor2_1 U28198 ( .ip1(\x[24][10] ), .ip2(n24370), .op(n24033) );
  not_ab_or_c_or_d U28199 ( .ip1(sig_in[11]), .ip2(n24035), .ip3(n24034), 
        .ip4(n24033), .op(n24036) );
  nor2_1 U28200 ( .ip1(n24037), .ip2(n24036), .op(n24313) );
  inv_1 U28201 ( .ip(n24313), .op(n24038) );
  nand2_1 U28202 ( .ip1(n24305), .ip2(n24038), .op(n24042) );
  and2_1 U28203 ( .ip1(n24235), .ip2(\x[24][13] ), .op(n24039) );
  or2_1 U28204 ( .ip1(\x[24][14] ), .ip2(n24039), .op(n24041) );
  or2_1 U28205 ( .ip1(n24230), .ip2(n24039), .op(n24040) );
  nand2_1 U28206 ( .ip1(n24041), .ip2(n24040), .op(n24304) );
  nand2_1 U28207 ( .ip1(\x[24][12] ), .ip2(n24079), .op(n24311) );
  nand3_1 U28208 ( .ip1(n24042), .ip2(n24304), .ip3(n24311), .op(n24089) );
  nor2_1 U28209 ( .ip1(\x[24][15] ), .ip2(n24090), .op(n24302) );
  nor2_1 U28210 ( .ip1(\x[25][15] ), .ip2(n24090), .op(n24080) );
  nor3_1 U28211 ( .ip1(\x[25][14] ), .ip2(n24080), .ip3(n24185), .op(n24088)
         );
  inv_1 U28212 ( .ip(\x[25][11] ), .op(n24078) );
  nor2_1 U28213 ( .ip1(\x[25][8] ), .ip2(n24100), .op(n24065) );
  nor2_1 U28214 ( .ip1(\x[25][9] ), .ip2(n24043), .op(n24066) );
  nor2_1 U28215 ( .ip1(\x[25][7] ), .ip2(n24044), .op(n24064) );
  and2_1 U28216 ( .ip1(n24461), .ip2(\x[25][7] ), .op(n24060) );
  nor3_1 U28217 ( .ip1(n24045), .ip2(\x[25][6] ), .ip3(n24060), .op(n24062) );
  nor2_1 U28218 ( .ip1(\x[25][5] ), .ip2(n24350), .op(n24055) );
  inv_1 U28219 ( .ip(\x[25][4] ), .op(n24046) );
  nor3_1 U28220 ( .ip1(sig_in[4]), .ip2(n24055), .ip3(n24046), .op(n24058) );
  and2_1 U28221 ( .ip1(n24335), .ip2(\x[25][2] ), .op(n24052) );
  nand2_1 U28222 ( .ip1(\x[25][1] ), .ip2(n20652), .op(n24050) );
  nand2_1 U28223 ( .ip1(\x[25][0] ), .ip2(n24143), .op(n24049) );
  nor2_1 U28224 ( .ip1(\x[25][2] ), .ip2(n24463), .op(n24048) );
  nor2_1 U28225 ( .ip1(\x[25][1] ), .ip2(n20652), .op(n24047) );
  not_ab_or_c_or_d U28226 ( .ip1(n24050), .ip2(n24049), .ip3(n24048), .ip4(
        n24047), .op(n24051) );
  not_ab_or_c_or_d U28227 ( .ip1(\x[25][3] ), .ip2(n22795), .ip3(n24052), 
        .ip4(n24051), .op(n24056) );
  nor2_1 U28228 ( .ip1(\x[25][3] ), .ip2(n22795), .op(n24054) );
  nor2_1 U28229 ( .ip1(\x[25][4] ), .ip2(n24256), .op(n24053) );
  nor4_1 U28230 ( .ip1(n24056), .ip2(n24055), .ip3(n24054), .ip4(n24053), .op(
        n24057) );
  ab_or_c_or_d U28231 ( .ip1(\x[25][5] ), .ip2(n24350), .ip3(n24058), .ip4(
        n24057), .op(n24059) );
  not_ab_or_c_or_d U28232 ( .ip1(\x[25][6] ), .ip2(n24045), .ip3(n24060), 
        .ip4(n24059), .op(n24061) );
  or2_1 U28233 ( .ip1(n24062), .ip2(n24061), .op(n24063) );
  nor4_1 U28234 ( .ip1(n24065), .ip2(n24066), .ip3(n24064), .ip4(n24063), .op(
        n24072) );
  nand2_1 U28235 ( .ip1(n24455), .ip2(\x[25][9] ), .op(n24070) );
  inv_1 U28236 ( .ip(n24066), .op(n24067) );
  nand3_1 U28237 ( .ip1(\x[25][8] ), .ip2(n23804), .ip3(n24067), .op(n24069)
         );
  nand2_1 U28238 ( .ip1(\x[25][11] ), .ip2(n24239), .op(n24068) );
  nand3_1 U28239 ( .ip1(n24070), .ip2(n24069), .ip3(n24068), .op(n24071) );
  not_ab_or_c_or_d U28240 ( .ip1(\x[25][10] ), .ip2(n24370), .ip3(n24072), 
        .ip4(n24071), .op(n24077) );
  inv_1 U28241 ( .ip(\x[25][12] ), .op(n24075) );
  not_ab_or_c_or_d U28242 ( .ip1(\x[25][11] ), .ip2(n24136), .ip3(\x[25][10] ), 
        .ip4(n23980), .op(n24074) );
  nor2_1 U28243 ( .ip1(\x[25][13] ), .ip2(n24376), .op(n24073) );
  ab_or_c_or_d U28244 ( .ip1(n17845), .ip2(n24075), .ip3(n24074), .ip4(n24073), 
        .op(n24076) );
  not_ab_or_c_or_d U28245 ( .ip1(sig_in[11]), .ip2(n24078), .ip3(n24077), 
        .ip4(n24076), .op(n24086) );
  nand2_1 U28246 ( .ip1(n24079), .ip2(\x[25][12] ), .op(n24084) );
  inv_1 U28247 ( .ip(n24080), .op(n24083) );
  nand2_1 U28248 ( .ip1(\x[25][13] ), .ip2(n24081), .op(n24082) );
  nand3_1 U28249 ( .ip1(n24084), .ip2(n24083), .ip3(n24082), .op(n24085) );
  not_ab_or_c_or_d U28250 ( .ip1(\x[25][14] ), .ip2(n24230), .ip3(n24086), 
        .ip4(n24085), .op(n24087) );
  ab_or_c_or_d U28251 ( .ip1(\x[25][15] ), .ip2(n24329), .ip3(n24088), .ip4(
        n24087), .op(n24287) );
  not_ab_or_c_or_d U28252 ( .ip1(n24301), .ip2(n24089), .ip3(n24302), .ip4(
        n24287), .op(n24709) );
  nand2_1 U28253 ( .ip1(\x[27][15] ), .ip2(n24329), .op(n24193) );
  and2_1 U28254 ( .ip1(n24332), .ip2(\x[27][13] ), .op(n24091) );
  nor2_1 U28255 ( .ip1(\x[27][15] ), .ip2(n24090), .op(n24288) );
  not_ab_or_c_or_d U28256 ( .ip1(\x[27][14] ), .ip2(n24230), .ip3(n24091), 
        .ip4(n24288), .op(n24295) );
  nand2_1 U28257 ( .ip1(\x[27][12] ), .ip2(n24233), .op(n24292) );
  nand2_1 U28258 ( .ip1(n24295), .ip2(n24292), .op(n24192) );
  nand2_1 U28259 ( .ip1(\x[27][9] ), .ip2(n24269), .op(n24094) );
  nor2_1 U28260 ( .ip1(\x[27][11] ), .ip2(n24456), .op(n24093) );
  nor2_1 U28261 ( .ip1(\x[27][10] ), .ip2(n24370), .op(n24092) );
  or2_1 U28262 ( .ip1(n24093), .ip2(n24092), .op(n24098) );
  or2_1 U28263 ( .ip1(n24094), .ip2(n24098), .op(n24097) );
  nand2_1 U28264 ( .ip1(\x[27][10] ), .ip2(n24370), .op(n24095) );
  or2_1 U28265 ( .ip1(n24095), .ip2(n24098), .op(n24096) );
  nand2_1 U28266 ( .ip1(n24097), .ip2(n24096), .op(n24135) );
  nor2_1 U28267 ( .ip1(n24164), .ip2(\x[27][9] ), .op(n24099) );
  nor2_1 U28268 ( .ip1(n24099), .ip2(n24098), .op(n24131) );
  inv_1 U28269 ( .ip(\x[27][7] ), .op(n24129) );
  nor2_1 U28270 ( .ip1(\x[27][8] ), .ip2(n24100), .op(n24128) );
  nor2_1 U28271 ( .ip1(\x[27][5] ), .ip2(n24350), .op(n24114) );
  inv_1 U28272 ( .ip(\x[27][4] ), .op(n24101) );
  nor3_1 U28273 ( .ip1(sig_in[4]), .ip2(n24114), .ip3(n24101), .op(n24117) );
  and2_1 U28274 ( .ip1(n24335), .ip2(\x[27][2] ), .op(n24111) );
  inv_1 U28275 ( .ip(\x[27][1] ), .op(n24103) );
  inv_1 U28276 ( .ip(\x[27][0] ), .op(n24102) );
  not_ab_or_c_or_d U28277 ( .ip1(n24464), .ip2(n24103), .ip3(sig_in[0]), .ip4(
        n24102), .op(n24104) );
  or2_1 U28278 ( .ip1(\x[27][1] ), .ip2(n24104), .op(n24106) );
  or2_1 U28279 ( .ip1(n21685), .ip2(n24104), .op(n24105) );
  nand2_1 U28280 ( .ip1(n24106), .ip2(n24105), .op(n24109) );
  nor2_1 U28281 ( .ip1(\x[27][2] ), .ip2(n24107), .op(n24108) );
  nor2_1 U28282 ( .ip1(n24109), .ip2(n24108), .op(n24110) );
  not_ab_or_c_or_d U28283 ( .ip1(\x[27][3] ), .ip2(n24342), .ip3(n24111), 
        .ip4(n24110), .op(n24115) );
  nor2_1 U28284 ( .ip1(\x[27][4] ), .ip2(n24256), .op(n24113) );
  nor2_1 U28285 ( .ip1(\x[27][3] ), .ip2(n22525), .op(n24112) );
  nor4_1 U28286 ( .ip1(n24115), .ip2(n24114), .ip3(n24113), .ip4(n24112), .op(
        n24116) );
  not_ab_or_c_or_d U28287 ( .ip1(\x[27][6] ), .ip2(n23770), .ip3(n24117), 
        .ip4(n24116), .op(n24118) );
  nor2_1 U28288 ( .ip1(\x[27][6] ), .ip2(n24355), .op(n24120) );
  or2_1 U28289 ( .ip1(n24118), .ip2(n24120), .op(n24123) );
  nand2_1 U28290 ( .ip1(\x[27][5] ), .ip2(n24119), .op(n24121) );
  or2_1 U28291 ( .ip1(n24121), .ip2(n24120), .op(n24122) );
  nand2_1 U28292 ( .ip1(n24123), .ip2(n24122), .op(n24124) );
  or2_1 U28293 ( .ip1(\x[27][7] ), .ip2(n24124), .op(n24126) );
  or2_1 U28294 ( .ip1(n24044), .ip2(n24124), .op(n24125) );
  nand2_1 U28295 ( .ip1(n24126), .ip2(n24125), .op(n24127) );
  not_ab_or_c_or_d U28296 ( .ip1(sig_in[7]), .ip2(n24129), .ip3(n24128), .ip4(
        n24127), .op(n24130) );
  nand2_1 U28297 ( .ip1(n24131), .ip2(n24130), .op(n24133) );
  nand3_1 U28298 ( .ip1(n24131), .ip2(n23804), .ip3(\x[27][8] ), .op(n24132)
         );
  nand2_1 U28299 ( .ip1(n24133), .ip2(n24132), .op(n24134) );
  not_ab_or_c_or_d U28300 ( .ip1(\x[27][11] ), .ip2(n24136), .ip3(n24135), 
        .ip4(n24134), .op(n24291) );
  nor2_1 U28301 ( .ip1(\x[27][13] ), .ip2(n24137), .op(n24139) );
  nor2_1 U28302 ( .ip1(\x[27][12] ), .ip2(n24450), .op(n24138) );
  nor2_1 U28303 ( .ip1(n24139), .ip2(n24138), .op(n24293) );
  inv_1 U28304 ( .ip(n24293), .op(n24141) );
  or2_1 U28305 ( .ip1(n24185), .ip2(\x[27][14] ), .op(n24140) );
  nand2_1 U28306 ( .ip1(n24140), .ip2(n24193), .op(n24289) );
  nor3_1 U28307 ( .ip1(n24291), .ip2(n24141), .ip3(n24289), .op(n24191) );
  nand2_1 U28308 ( .ip1(\x[28][8] ), .ip2(n23804), .op(n24163) );
  nor2_1 U28309 ( .ip1(n24142), .ip2(\x[28][7] ), .op(n24161) );
  inv_1 U28310 ( .ip(\x[28][5] ), .op(n24157) );
  nor2_1 U28311 ( .ip1(sig_in[5]), .ip2(n24157), .op(n24154) );
  inv_1 U28312 ( .ip(\x[28][3] ), .op(n24152) );
  and2_1 U28313 ( .ip1(n24335), .ip2(\x[28][2] ), .op(n24149) );
  nand2_1 U28314 ( .ip1(\x[28][1] ), .ip2(n20652), .op(n24147) );
  nand2_1 U28315 ( .ip1(\x[28][0] ), .ip2(n24143), .op(n24146) );
  nor2_1 U28316 ( .ip1(\x[28][2] ), .ip2(n24463), .op(n24145) );
  nor2_1 U28317 ( .ip1(\x[28][1] ), .ip2(n20652), .op(n24144) );
  not_ab_or_c_or_d U28318 ( .ip1(n24147), .ip2(n24146), .ip3(n24145), .ip4(
        n24144), .op(n24148) );
  not_ab_or_c_or_d U28319 ( .ip1(\x[28][3] ), .ip2(n24476), .ip3(n24149), 
        .ip4(n24148), .op(n24151) );
  nor2_1 U28320 ( .ip1(\x[28][4] ), .ip2(n24256), .op(n24150) );
  not_ab_or_c_or_d U28321 ( .ip1(sig_in[3]), .ip2(n24152), .ip3(n24151), .ip4(
        n24150), .op(n24153) );
  not_ab_or_c_or_d U28322 ( .ip1(\x[28][4] ), .ip2(n24256), .ip3(n24154), 
        .ip4(n24153), .op(n24156) );
  nor2_1 U28323 ( .ip1(\x[28][6] ), .ip2(n24355), .op(n24155) );
  not_ab_or_c_or_d U28324 ( .ip1(n22833), .ip2(n24157), .ip3(n24156), .ip4(
        n24155), .op(n24159) );
  and2_1 U28325 ( .ip1(n23509), .ip2(\x[28][6] ), .op(n24158) );
  not_ab_or_c_or_d U28326 ( .ip1(\x[28][7] ), .ip2(n24492), .ip3(n24159), 
        .ip4(n24158), .op(n24160) );
  nor2_1 U28327 ( .ip1(n24161), .ip2(n24160), .op(n24203) );
  inv_1 U28328 ( .ip(n24203), .op(n24162) );
  nand2_1 U28329 ( .ip1(n24163), .ip2(n24162), .op(n24167) );
  nor2_1 U28330 ( .ip1(\x[28][9] ), .ip2(n24164), .op(n24195) );
  or2_1 U28331 ( .ip1(sig_in[8]), .ip2(n24195), .op(n24166) );
  inv_1 U28332 ( .ip(\x[28][8] ), .op(n24196) );
  or2_1 U28333 ( .ip1(n24196), .ip2(n24195), .op(n24165) );
  nand2_1 U28334 ( .ip1(n24166), .ip2(n24165), .op(n24201) );
  nand2_1 U28335 ( .ip1(n24167), .ip2(n24201), .op(n24169) );
  and2_1 U28336 ( .ip1(n24451), .ip2(\x[28][10] ), .op(n24168) );
  and2_1 U28337 ( .ip1(n24239), .ip2(\x[28][11] ), .op(n24172) );
  not_ab_or_c_or_d U28338 ( .ip1(\x[28][9] ), .ip2(n24455), .ip3(n24168), 
        .ip4(n24172), .op(n24198) );
  nand2_1 U28339 ( .ip1(n24169), .ip2(n24198), .op(n24173) );
  nor2_1 U28340 ( .ip1(\x[28][11] ), .ip2(n21793), .op(n24171) );
  nor2_1 U28341 ( .ip1(\x[28][10] ), .ip2(n24457), .op(n24170) );
  nor2_1 U28342 ( .ip1(n24171), .ip2(n24170), .op(n24202) );
  or2_1 U28343 ( .ip1(n24172), .ip2(n24202), .op(n24200) );
  nand2_1 U28344 ( .ip1(n24173), .ip2(n24200), .op(n24174) );
  nand2_1 U28345 ( .ip1(\x[28][12] ), .ip2(n24449), .op(n24214) );
  nand2_1 U28346 ( .ip1(n24174), .ip2(n24214), .op(n24179) );
  nor2_1 U28347 ( .ip1(\x[28][13] ), .ip2(n24376), .op(n24175) );
  or2_1 U28348 ( .ip1(sig_in[12]), .ip2(n24175), .op(n24178) );
  inv_1 U28349 ( .ip(\x[28][12] ), .op(n24176) );
  or2_1 U28350 ( .ip1(n24176), .ip2(n24175), .op(n24177) );
  nand2_1 U28351 ( .ip1(n24178), .ip2(n24177), .op(n24204) );
  nand2_1 U28352 ( .ip1(n24179), .ip2(n24204), .op(n24183) );
  nor2_1 U28353 ( .ip1(\x[28][15] ), .ip2(n24180), .op(n24184) );
  nand2_1 U28354 ( .ip1(n24235), .ip2(\x[28][13] ), .op(n24213) );
  inv_1 U28355 ( .ip(n24213), .op(n24181) );
  not_ab_or_c_or_d U28356 ( .ip1(\x[28][14] ), .ip2(n24382), .ip3(n24184), 
        .ip4(n24181), .op(n24182) );
  nand2_1 U28357 ( .ip1(n24183), .ip2(n24182), .op(n24189) );
  inv_1 U28358 ( .ip(n24184), .op(n24209) );
  or2_1 U28359 ( .ip1(n24185), .ip2(\x[28][14] ), .op(n24187) );
  nand2_1 U28360 ( .ip1(\x[28][15] ), .ip2(n24186), .op(n24210) );
  nand2_1 U28361 ( .ip1(n24187), .ip2(n24210), .op(n24212) );
  nand2_1 U28362 ( .ip1(n24209), .ip2(n24212), .op(n24188) );
  nand2_1 U28363 ( .ip1(n24189), .ip2(n24188), .op(n24190) );
  not_ab_or_c_or_d U28364 ( .ip1(n24193), .ip2(n24192), .ip3(n24191), .ip4(
        n24190), .op(n27398) );
  inv_1 U28365 ( .ip(n24194), .op(n24225) );
  or3_1 U28366 ( .ip1(n23779), .ip2(n24196), .ip3(n24195), .op(n24197) );
  nand2_1 U28367 ( .ip1(n24198), .ip2(n24197), .op(n24199) );
  nand2_1 U28368 ( .ip1(n24200), .ip2(n24199), .op(n24207) );
  nand3_1 U28369 ( .ip1(n24203), .ip2(n24202), .ip3(n24201), .op(n24206) );
  inv_1 U28370 ( .ip(n24204), .op(n24205) );
  not_ab_or_c_or_d U28371 ( .ip1(n24207), .ip2(n24206), .ip3(n24205), .ip4(
        n24212), .op(n24224) );
  nand2_1 U28372 ( .ip1(\x[28][14] ), .ip2(n24327), .op(n24208) );
  nand2_1 U28373 ( .ip1(n24209), .ip2(n24208), .op(n24211) );
  nand2_1 U28374 ( .ip1(n24211), .ip2(n24210), .op(n24221) );
  inv_1 U28375 ( .ip(n24212), .op(n24216) );
  nand2_1 U28376 ( .ip1(n24214), .ip2(n24213), .op(n24215) );
  nand2_1 U28377 ( .ip1(n24216), .ip2(n24215), .op(n24220) );
  or2_1 U28378 ( .ip1(n24218), .ip2(n24217), .op(n24219) );
  nand4_1 U28379 ( .ip1(n24222), .ip2(n24221), .ip3(n24220), .ip4(n24219), 
        .op(n24223) );
  not_ab_or_c_or_d U28380 ( .ip1(n24226), .ip2(n24225), .ip3(n24224), .ip4(
        n24223), .op(n27400) );
  nor2_1 U28381 ( .ip1(n27398), .ip2(n27400), .op(n24704) );
  inv_1 U28382 ( .ip(\x[26][15] ), .op(n24229) );
  nor2_1 U28383 ( .ip1(n24229), .ip2(sig_in[15]), .op(n24228) );
  not_ab_or_c_or_d U28384 ( .ip1(sig_in[15]), .ip2(n24229), .ip3(\x[26][14] ), 
        .ip4(n24327), .op(n24227) );
  or2_1 U28385 ( .ip1(n24228), .ip2(n24227), .op(n24286) );
  nand2_1 U28386 ( .ip1(sig_in[15]), .ip2(n24229), .op(n24232) );
  nand2_1 U28387 ( .ip1(\x[26][14] ), .ip2(n24230), .op(n24231) );
  nand2_1 U28388 ( .ip1(n24232), .ip2(n24231), .op(n24234) );
  nor3_1 U28389 ( .ip1(\x[26][13] ), .ip2(n24235), .ip3(n24234), .op(n24285)
         );
  or2_1 U28390 ( .ip1(n24233), .ip2(\x[26][12] ), .op(n24238) );
  inv_1 U28391 ( .ip(n24234), .op(n24237) );
  nand2_1 U28392 ( .ip1(\x[26][13] ), .ip2(n24235), .op(n24236) );
  nand2_1 U28393 ( .ip1(n24237), .ip2(n24236), .op(n24280) );
  or2_1 U28394 ( .ip1(n24238), .ip2(n24280), .op(n24283) );
  nand2_1 U28395 ( .ip1(\x[26][11] ), .ip2(n24239), .op(n24279) );
  nor2_1 U28396 ( .ip1(\x[26][10] ), .ip2(n24457), .op(n24240) );
  or2_1 U28397 ( .ip1(sig_in[11]), .ip2(n24240), .op(n24243) );
  inv_1 U28398 ( .ip(\x[26][11] ), .op(n24241) );
  or2_1 U28399 ( .ip1(n24241), .ip2(n24240), .op(n24242) );
  nand2_1 U28400 ( .ip1(n24243), .ip2(n24242), .op(n24276) );
  nand2_1 U28401 ( .ip1(\x[26][10] ), .ip2(n24370), .op(n24274) );
  inv_1 U28402 ( .ip(\x[26][7] ), .op(n24265) );
  nor2_1 U28403 ( .ip1(n17732), .ip2(n24265), .op(n24262) );
  inv_1 U28404 ( .ip(\x[26][3] ), .op(n24250) );
  nor2_1 U28405 ( .ip1(\x[26][2] ), .ip2(n24463), .op(n24249) );
  inv_1 U28406 ( .ip(\x[26][1] ), .op(n24245) );
  nor2_1 U28407 ( .ip1(sig_in[1]), .ip2(n24245), .op(n24247) );
  inv_1 U28408 ( .ip(\x[26][0] ), .op(n24244) );
  not_ab_or_c_or_d U28409 ( .ip1(n24467), .ip2(n24245), .ip3(sig_in[0]), .ip4(
        n24244), .op(n24246) );
  not_ab_or_c_or_d U28410 ( .ip1(\x[26][2] ), .ip2(n24470), .ip3(n24247), 
        .ip4(n24246), .op(n24248) );
  not_ab_or_c_or_d U28411 ( .ip1(n24251), .ip2(n24250), .ip3(n24249), .ip4(
        n24248), .op(n24255) );
  nand2_1 U28412 ( .ip1(\x[26][5] ), .ip2(n24350), .op(n24253) );
  nand2_1 U28413 ( .ip1(\x[26][4] ), .ip2(n24347), .op(n24252) );
  nand2_1 U28414 ( .ip1(n24253), .ip2(n24252), .op(n24254) );
  not_ab_or_c_or_d U28415 ( .ip1(\x[26][3] ), .ip2(n24342), .ip3(n24255), 
        .ip4(n24254), .op(n24260) );
  nor2_1 U28416 ( .ip1(\x[26][5] ), .ip2(n24350), .op(n24259) );
  nor2_1 U28417 ( .ip1(\x[26][6] ), .ip2(n24355), .op(n24258) );
  not_ab_or_c_or_d U28418 ( .ip1(\x[26][5] ), .ip2(n24482), .ip3(\x[26][4] ), 
        .ip4(n24256), .op(n24257) );
  nor4_1 U28419 ( .ip1(n24260), .ip2(n24259), .ip3(n24258), .ip4(n24257), .op(
        n24261) );
  not_ab_or_c_or_d U28420 ( .ip1(\x[26][6] ), .ip2(n23770), .ip3(n24262), 
        .ip4(n24261), .op(n24264) );
  nor2_1 U28421 ( .ip1(\x[26][8] ), .ip2(n24358), .op(n24263) );
  not_ab_or_c_or_d U28422 ( .ip1(sig_in[7]), .ip2(n24265), .ip3(n24264), .ip4(
        n24263), .op(n24266) );
  or2_1 U28423 ( .ip1(\x[26][8] ), .ip2(n24266), .op(n24268) );
  or2_1 U28424 ( .ip1(n24491), .ip2(n24266), .op(n24267) );
  nand2_1 U28425 ( .ip1(n24268), .ip2(n24267), .op(n24271) );
  nor2_1 U28426 ( .ip1(\x[26][9] ), .ip2(n24269), .op(n24270) );
  or2_1 U28427 ( .ip1(n24271), .ip2(n24270), .op(n24273) );
  nand2_1 U28428 ( .ip1(\x[26][9] ), .ip2(n23981), .op(n24272) );
  nand3_1 U28429 ( .ip1(n24274), .ip2(n24273), .ip3(n24272), .op(n24275) );
  nand2_1 U28430 ( .ip1(n24276), .ip2(n24275), .op(n24278) );
  nand2_1 U28431 ( .ip1(\x[26][12] ), .ip2(n24450), .op(n24277) );
  nand3_1 U28432 ( .ip1(n24279), .ip2(n24278), .ip3(n24277), .op(n24281) );
  or2_1 U28433 ( .ip1(n24281), .ip2(n24280), .op(n24282) );
  nand2_1 U28434 ( .ip1(n24283), .ip2(n24282), .op(n24284) );
  nor3_1 U28435 ( .ip1(n24286), .ip2(n24285), .ip3(n24284), .op(n24297) );
  nand2_1 U28436 ( .ip1(n24297), .ip2(n24287), .op(n24705) );
  inv_1 U28437 ( .ip(n24288), .op(n24290) );
  nand2_1 U28438 ( .ip1(n24290), .ip2(n24289), .op(n24300) );
  nand2_1 U28439 ( .ip1(n24292), .ip2(n24291), .op(n24294) );
  nand2_1 U28440 ( .ip1(n24294), .ip2(n24293), .op(n24296) );
  nand2_1 U28441 ( .ip1(n24296), .ip2(n24295), .op(n24299) );
  inv_1 U28442 ( .ip(n24297), .op(n24298) );
  nand3_1 U28443 ( .ip1(n24300), .ip2(n24299), .ip3(n24298), .op(n24715) );
  nand3_1 U28444 ( .ip1(n24704), .ip2(n24705), .ip3(n24715), .op(n24710) );
  nor2_1 U28445 ( .ip1(n24709), .ip2(n24710), .op(n24712) );
  nor2_1 U28446 ( .ip1(n24302), .ip2(n24301), .op(n24307) );
  inv_1 U28447 ( .ip(n24302), .op(n24303) );
  nand2_1 U28448 ( .ip1(n24304), .ip2(n24303), .op(n24310) );
  nor2_1 U28449 ( .ip1(n24305), .ip2(n24310), .op(n24306) );
  not_ab_or_c_or_d U28450 ( .ip1(n24309), .ip2(n24308), .ip3(n24307), .ip4(
        n24306), .op(n24319) );
  inv_1 U28451 ( .ip(n24310), .op(n24312) );
  nand3_1 U28452 ( .ip1(n24313), .ip2(n24312), .ip3(n24311), .op(n24318) );
  nand3_1 U28453 ( .ip1(n24316), .ip2(n24315), .ip3(n24314), .op(n24317) );
  nand3_1 U28454 ( .ip1(n24319), .ip2(n24318), .ip3(n24317), .op(n24714) );
  nand2_1 U28455 ( .ip1(n24712), .ip2(n24714), .op(n24794) );
  nor2_1 U28456 ( .ip1(n24793), .ip2(n24794), .op(n24777) );
  inv_1 U28457 ( .ip(n24320), .op(n24321) );
  nand2_1 U28458 ( .ip1(n24322), .ip2(n24321), .op(n24324) );
  nand2_1 U28459 ( .ip1(n24324), .ip2(n24323), .op(n24326) );
  nand2_1 U28460 ( .ip1(n24326), .ip2(n24325), .op(n24387) );
  nor2_1 U28461 ( .ip1(\x[21][14] ), .ip2(n24327), .op(n24328) );
  or2_1 U28462 ( .ip1(\x[21][15] ), .ip2(n24328), .op(n24331) );
  or2_1 U28463 ( .ip1(n24329), .ip2(n24328), .op(n24330) );
  nand2_1 U28464 ( .ip1(n24331), .ip2(n24330), .op(n24393) );
  and2_1 U28465 ( .ip1(n24332), .ip2(\x[21][13] ), .op(n24381) );
  inv_1 U28466 ( .ip(\x[21][12] ), .op(n24379) );
  inv_1 U28467 ( .ip(\x[21][9] ), .op(n24334) );
  nor2_1 U28468 ( .ip1(\x[21][10] ), .ip2(n24457), .op(n24333) );
  nor2_1 U28469 ( .ip1(\x[21][11] ), .ip2(n24456), .op(n24368) );
  not_ab_or_c_or_d U28470 ( .ip1(sig_in[9]), .ip2(n24334), .ip3(n24333), .ip4(
        n24368), .op(n24367) );
  and2_1 U28471 ( .ip1(n24355), .ip2(\x[21][6] ), .op(n24354) );
  inv_1 U28472 ( .ip(\x[21][3] ), .op(n24345) );
  and2_1 U28473 ( .ip1(n24335), .ip2(\x[21][2] ), .op(n24341) );
  nand2_1 U28474 ( .ip1(\x[21][1] ), .ip2(n21685), .op(n24339) );
  nand2_1 U28475 ( .ip1(\x[21][0] ), .ip2(n24143), .op(n24338) );
  nor2_1 U28476 ( .ip1(\x[21][2] ), .ip2(n24463), .op(n24337) );
  nor2_1 U28477 ( .ip1(\x[21][1] ), .ip2(n21685), .op(n24336) );
  not_ab_or_c_or_d U28478 ( .ip1(n24339), .ip2(n24338), .ip3(n24337), .ip4(
        n24336), .op(n24340) );
  not_ab_or_c_or_d U28479 ( .ip1(\x[21][3] ), .ip2(n24342), .ip3(n24341), 
        .ip4(n24340), .op(n24344) );
  nor2_1 U28480 ( .ip1(\x[21][4] ), .ip2(n23721), .op(n24343) );
  not_ab_or_c_or_d U28481 ( .ip1(sig_in[3]), .ip2(n24345), .ip3(n24344), .ip4(
        n24343), .op(n24346) );
  or2_1 U28482 ( .ip1(\x[21][4] ), .ip2(n24346), .op(n24349) );
  or2_1 U28483 ( .ip1(n24347), .ip2(n24346), .op(n24348) );
  nand2_1 U28484 ( .ip1(n24349), .ip2(n24348), .op(n24352) );
  nor2_1 U28485 ( .ip1(\x[21][5] ), .ip2(n24350), .op(n24351) );
  nor2_1 U28486 ( .ip1(n24352), .ip2(n24351), .op(n24353) );
  not_ab_or_c_or_d U28487 ( .ip1(\x[21][5] ), .ip2(n24482), .ip3(n24354), 
        .ip4(n24353), .op(n24357) );
  nor2_1 U28488 ( .ip1(\x[21][6] ), .ip2(n24355), .op(n24356) );
  nor2_1 U28489 ( .ip1(n24357), .ip2(n24356), .op(n24359) );
  nand2_1 U28490 ( .ip1(n24359), .ip2(\x[21][7] ), .op(n24362) );
  nor2_1 U28491 ( .ip1(\x[21][8] ), .ip2(n24358), .op(n24361) );
  nor2_1 U28492 ( .ip1(n24359), .ip2(\x[21][7] ), .op(n24360) );
  ab_or_c_or_d U28493 ( .ip1(n17732), .ip2(n24362), .ip3(n24361), .ip4(n24360), 
        .op(n24365) );
  nand2_1 U28494 ( .ip1(\x[21][9] ), .ip2(n24043), .op(n24364) );
  nand2_1 U28495 ( .ip1(\x[21][8] ), .ip2(n24491), .op(n24363) );
  nand3_1 U28496 ( .ip1(n24365), .ip2(n24364), .ip3(n24363), .op(n24366) );
  nand2_1 U28497 ( .ip1(n24367), .ip2(n24366), .op(n24375) );
  inv_1 U28498 ( .ip(n24368), .op(n24369) );
  nand3_1 U28499 ( .ip1(\x[21][10] ), .ip2(n24370), .ip3(n24369), .op(n24374)
         );
  nand2_1 U28500 ( .ip1(\x[21][12] ), .ip2(n24450), .op(n24373) );
  nand2_1 U28501 ( .ip1(\x[21][11] ), .ip2(n24371), .op(n24372) );
  and4_1 U28502 ( .ip1(n24375), .ip2(n24374), .ip3(n24373), .ip4(n24372), .op(
        n24378) );
  nor2_1 U28503 ( .ip1(\x[21][13] ), .ip2(n24376), .op(n24377) );
  not_ab_or_c_or_d U28504 ( .ip1(sig_in[12]), .ip2(n24379), .ip3(n24378), 
        .ip4(n24377), .op(n24380) );
  not_ab_or_c_or_d U28505 ( .ip1(\x[21][14] ), .ip2(n24382), .ip3(n24381), 
        .ip4(n24380), .op(n24397) );
  inv_1 U28506 ( .ip(n24397), .op(n24383) );
  nand2_1 U28507 ( .ip1(n24393), .ip2(n24383), .op(n24385) );
  nor2_1 U28508 ( .ip1(n24384), .ip2(\x[21][15] ), .op(n24392) );
  inv_1 U28509 ( .ip(n24392), .op(n24396) );
  nand4_1 U28510 ( .ip1(n24387), .ip2(n24386), .ip3(n24385), .ip4(n24396), 
        .op(n24778) );
  nand2_1 U28511 ( .ip1(n24389), .ip2(n24388), .op(n24391) );
  nand2_1 U28512 ( .ip1(n24391), .ip2(n24390), .op(n24404) );
  nor2_1 U28513 ( .ip1(n24393), .ip2(n24392), .op(n24394) );
  not_ab_or_c_or_d U28514 ( .ip1(n24397), .ip2(n24396), .ip3(n24395), .ip4(
        n24394), .op(n24403) );
  inv_1 U28515 ( .ip(n24398), .op(n24399) );
  nand3_1 U28516 ( .ip1(n24401), .ip2(n24400), .ip3(n24399), .op(n24402) );
  nand3_1 U28517 ( .ip1(n24404), .ip2(n24403), .ip3(n24402), .op(n24779) );
  nand3_1 U28518 ( .ip1(n24777), .ip2(n24778), .ip3(n24779), .op(n24791) );
  nor2_1 U28519 ( .ip1(n24790), .ip2(n24791), .op(n24774) );
  nand2_1 U28520 ( .ip1(n24406), .ip2(n24405), .op(n24408) );
  nand2_1 U28521 ( .ip1(n24408), .ip2(n24407), .op(n24425) );
  inv_1 U28522 ( .ip(n24409), .op(n24417) );
  and2_1 U28523 ( .ip1(n24411), .ip2(n24410), .op(n24416) );
  inv_1 U28524 ( .ip(n24412), .op(n24413) );
  nor2_1 U28525 ( .ip1(n24414), .ip2(n24413), .op(n24415) );
  not_ab_or_c_or_d U28526 ( .ip1(n24418), .ip2(n24417), .ip3(n24416), .ip4(
        n24415), .op(n24424) );
  inv_1 U28527 ( .ip(n24419), .op(n24420) );
  or3_1 U28528 ( .ip1(n24422), .ip2(n24421), .ip3(n24420), .op(n24423) );
  nand3_1 U28529 ( .ip1(n24425), .ip2(n24424), .ip3(n24423), .op(n24776) );
  nand2_1 U28530 ( .ip1(n24774), .ip2(n24776), .op(n24703) );
  nor2_1 U28531 ( .ip1(n24701), .ip2(n24703), .op(n24781) );
  inv_1 U28532 ( .ip(n24426), .op(n24427) );
  nor2_1 U28533 ( .ip1(n24427), .ip2(n24429), .op(n24443) );
  inv_1 U28534 ( .ip(n24428), .op(n24432) );
  nor3_1 U28535 ( .ip1(\x[17][14] ), .ip2(n24429), .ip3(n24382), .op(n24430)
         );
  not_ab_or_c_or_d U28536 ( .ip1(n24443), .ip2(n24432), .ip3(n24431), .ip4(
        n24430), .op(n24448) );
  inv_1 U28537 ( .ip(n24433), .op(n24440) );
  nand2_1 U28538 ( .ip1(n24435), .ip2(n24434), .op(n24438) );
  nand3_1 U28539 ( .ip1(n24438), .ip2(n24437), .ip3(n24436), .op(n24439) );
  nand2_1 U28540 ( .ip1(n24440), .ip2(n24439), .op(n24447) );
  inv_1 U28541 ( .ip(n24441), .op(n24442) );
  nand3_1 U28542 ( .ip1(n24444), .ip2(n24443), .ip3(n24442), .op(n24445) );
  nand4_1 U28543 ( .ip1(n24448), .ip2(n24447), .ip3(n24446), .ip4(n24445), 
        .op(n24782) );
  nand2_1 U28544 ( .ip1(n24781), .ip2(n24782), .op(n24724) );
  nor2_1 U28545 ( .ip1(n24722), .ip2(n24724), .op(n24772) );
  inv_1 U28546 ( .ip(\x[0][13] ), .op(n24505) );
  nor2_1 U28547 ( .ip1(n24505), .ip2(sig_in[13]), .op(n24507) );
  nor2_1 U28548 ( .ip1(\x[0][12] ), .ip2(n24449), .op(n24504) );
  and2_1 U28549 ( .ip1(n24450), .ip2(\x[0][12] ), .op(n24502) );
  and2_1 U28550 ( .ip1(n24451), .ip2(\x[0][10] ), .op(n24454) );
  nor2_1 U28551 ( .ip1(\x[0][9] ), .ip2(n24269), .op(n24494) );
  inv_1 U28552 ( .ip(\x[0][8] ), .op(n24452) );
  nor3_1 U28553 ( .ip1(sig_in[8]), .ip2(n24494), .ip3(n24452), .op(n24453) );
  not_ab_or_c_or_d U28554 ( .ip1(\x[0][9] ), .ip2(n24455), .ip3(n24454), .ip4(
        n24453), .op(n24460) );
  nor2_1 U28555 ( .ip1(\x[0][11] ), .ip2(n24456), .op(n24459) );
  nor2_1 U28556 ( .ip1(\x[0][10] ), .ip2(n24457), .op(n24458) );
  or2_1 U28557 ( .ip1(n24459), .ip2(n24458), .op(n24497) );
  or2_1 U28558 ( .ip1(n24460), .ip2(n24497), .op(n24500) );
  and2_1 U28559 ( .ip1(n24461), .ip2(\x[0][7] ), .op(n24490) );
  inv_1 U28560 ( .ip(\x[0][5] ), .op(n24488) );
  inv_1 U28561 ( .ip(\x[0][4] ), .op(n24478) );
  nor2_1 U28562 ( .ip1(n24462), .ip2(n24478), .op(n24475) );
  inv_1 U28563 ( .ip(\x[0][3] ), .op(n24473) );
  nor2_1 U28564 ( .ip1(\x[0][2] ), .ip2(n24463), .op(n24472) );
  inv_1 U28565 ( .ip(\x[0][1] ), .op(n24466) );
  nor2_1 U28566 ( .ip1(n24464), .ip2(n24466), .op(n24469) );
  inv_1 U28567 ( .ip(\x[0][0] ), .op(n24465) );
  not_ab_or_c_or_d U28568 ( .ip1(n24467), .ip2(n24466), .ip3(sig_in[0]), .ip4(
        n24465), .op(n24468) );
  not_ab_or_c_or_d U28569 ( .ip1(\x[0][2] ), .ip2(n24470), .ip3(n24469), .ip4(
        n24468), .op(n24471) );
  not_ab_or_c_or_d U28570 ( .ip1(n24251), .ip2(n24473), .ip3(n24472), .ip4(
        n24471), .op(n24474) );
  not_ab_or_c_or_d U28571 ( .ip1(\x[0][3] ), .ip2(n24476), .ip3(n24475), .ip4(
        n24474), .op(n24477) );
  or2_1 U28572 ( .ip1(sig_in[4]), .ip2(n24477), .op(n24480) );
  or2_1 U28573 ( .ip1(n24478), .ip2(n24477), .op(n24479) );
  nand2_1 U28574 ( .ip1(n24480), .ip2(n24479), .op(n24481) );
  or2_1 U28575 ( .ip1(\x[0][5] ), .ip2(n24481), .op(n24484) );
  or2_1 U28576 ( .ip1(n24482), .ip2(n24481), .op(n24483) );
  nand2_1 U28577 ( .ip1(n24484), .ip2(n24483), .op(n24487) );
  nor2_1 U28578 ( .ip1(\x[0][6] ), .ip2(n24485), .op(n24486) );
  not_ab_or_c_or_d U28579 ( .ip1(sig_in[5]), .ip2(n24488), .ip3(n24487), .ip4(
        n24486), .op(n24489) );
  not_ab_or_c_or_d U28580 ( .ip1(\x[0][6] ), .ip2(n23509), .ip3(n24490), .ip4(
        n24489), .op(n24496) );
  nor2_1 U28581 ( .ip1(\x[0][8] ), .ip2(n24491), .op(n24495) );
  nor2_1 U28582 ( .ip1(\x[0][7] ), .ip2(n24492), .op(n24493) );
  or4_1 U28583 ( .ip1(n24496), .ip2(n24495), .ip3(n24494), .ip4(n24493), .op(
        n24498) );
  or2_1 U28584 ( .ip1(n24498), .ip2(n24497), .op(n24499) );
  nand2_1 U28585 ( .ip1(n24500), .ip2(n24499), .op(n24501) );
  not_ab_or_c_or_d U28586 ( .ip1(\x[0][11] ), .ip2(n24371), .ip3(n24502), 
        .ip4(n24501), .op(n24503) );
  not_ab_or_c_or_d U28587 ( .ip1(sig_in[13]), .ip2(n24505), .ip3(n24504), 
        .ip4(n24503), .op(n24506) );
  or2_1 U28588 ( .ip1(n24507), .ip2(n24506), .op(n24508) );
  nand2_1 U28589 ( .ip1(\x[0][14] ), .ip2(n24508), .op(n24511) );
  inv_1 U28590 ( .ip(\x[0][15] ), .op(n24512) );
  nor2_1 U28591 ( .ip1(sig_in[15]), .ip2(n24512), .op(n24510) );
  nor2_1 U28592 ( .ip1(\x[0][14] ), .ip2(n24508), .op(n24509) );
  ab_or_c_or_d U28593 ( .ip1(sig_in[14]), .ip2(n24511), .ip3(n24510), .ip4(
        n24509), .op(n24516) );
  nand2_1 U28594 ( .ip1(sig_in[15]), .ip2(n24512), .op(n24513) );
  nand4_1 U28595 ( .ip1(n24516), .ip2(n24515), .ip3(n24514), .ip4(n24513), 
        .op(n24517) );
  and4_1 U28596 ( .ip1(n27436), .ip2(n24518), .ip3(n24772), .ip4(n24517), .op(
        n24519) );
  nand4_1 U28597 ( .ip1(n27533), .ip2(n27567), .ip3(n27288), .ip4(n24519), 
        .op(n24967) );
  nand2_1 U28598 ( .ip1(n26295), .ip2(n24967), .op(n24520) );
  nor2_1 U28599 ( .ip1(n24521), .ip2(n24520), .op(n27589) );
  inv_1 U28600 ( .ip(n24522), .op(n24523) );
  nand2_1 U28601 ( .ip1(n24524), .ip2(n24523), .op(n25965) );
  nor2_1 U28602 ( .ip1(n27371), .ip2(n25965), .op(n27581) );
  inv_1 U28603 ( .ip(n24525), .op(n27364) );
  nor2_1 U28604 ( .ip1(n27364), .ip2(n27367), .op(n27156) );
  inv_1 U28605 ( .ip(n24526), .op(n24527) );
  nor2_1 U28606 ( .ip1(n24528), .ip2(n24527), .op(n27363) );
  inv_1 U28607 ( .ip(n24529), .op(n24531) );
  nor2_1 U28608 ( .ip1(n24531), .ip2(n24530), .op(n27349) );
  inv_1 U28609 ( .ip(n24532), .op(n24533) );
  nor2_1 U28610 ( .ip1(n24534), .ip2(n24533), .op(n27333) );
  nand2_1 U28611 ( .ip1(n27333), .ip2(\LUT[95][0] ), .op(n24541) );
  inv_1 U28612 ( .ip(n24535), .op(n24537) );
  nor2_1 U28613 ( .ip1(n24537), .ip2(n24536), .op(n27334) );
  nand2_1 U28614 ( .ip1(n27334), .ip2(\LUT[94][0] ), .op(n24540) );
  nand2_1 U28615 ( .ip1(n27335), .ip2(\LUT[98][0] ), .op(n24539) );
  nand2_1 U28616 ( .ip1(n27336), .ip2(\LUT[97][0] ), .op(n24538) );
  nand4_1 U28617 ( .ip1(n24541), .ip2(n24540), .ip3(n24539), .ip4(n24538), 
        .op(n24555) );
  inv_1 U28618 ( .ip(n24542), .op(n24543) );
  nor2_1 U28619 ( .ip1(n24544), .ip2(n24543), .op(n27341) );
  nand2_1 U28620 ( .ip1(n27341), .ip2(\LUT[93][0] ), .op(n24553) );
  inv_1 U28621 ( .ip(n24545), .op(n24547) );
  nor2_1 U28622 ( .ip1(n24547), .ip2(n24546), .op(n27342) );
  nand2_1 U28623 ( .ip1(n27342), .ip2(\LUT[92][0] ), .op(n24552) );
  inv_1 U28624 ( .ip(n24548), .op(n24550) );
  nor2_1 U28625 ( .ip1(n24550), .ip2(n24549), .op(n27343) );
  nand2_1 U28626 ( .ip1(n27343), .ip2(\LUT[91][0] ), .op(n24551) );
  nand3_1 U28627 ( .ip1(n24553), .ip2(n24552), .ip3(n24551), .op(n24554) );
  not_ab_or_c_or_d U28628 ( .ip1(n27349), .ip2(\LUT[96][0] ), .ip3(n24555), 
        .ip4(n24554), .op(n24568) );
  inv_1 U28629 ( .ip(n24556), .op(n24557) );
  nor2_1 U28630 ( .ip1(n24558), .ip2(n24557), .op(n27350) );
  nand2_1 U28631 ( .ip1(n27350), .ip2(\LUT[89][0] ), .op(n24567) );
  inv_1 U28632 ( .ip(n24559), .op(n24560) );
  nor2_1 U28633 ( .ip1(n24561), .ip2(n24560), .op(n27351) );
  nand2_1 U28634 ( .ip1(n27351), .ip2(\LUT[90][0] ), .op(n24566) );
  inv_1 U28635 ( .ip(n24562), .op(n24564) );
  nor2_1 U28636 ( .ip1(n24564), .ip2(n24563), .op(n27352) );
  nand2_1 U28637 ( .ip1(n27352), .ip2(\LUT[88][0] ), .op(n24565) );
  nand4_1 U28638 ( .ip1(n24568), .ip2(n24567), .ip3(n24566), .ip4(n24565), 
        .op(n24578) );
  inv_1 U28639 ( .ip(n24569), .op(n24570) );
  nor2_1 U28640 ( .ip1(n24571), .ip2(n24570), .op(n27357) );
  nand2_1 U28641 ( .ip1(\LUT[85][0] ), .ip2(n27357), .op(n24576) );
  inv_1 U28642 ( .ip(n24572), .op(n24574) );
  nor2_1 U28643 ( .ip1(n24574), .ip2(n24573), .op(n27358) );
  nand2_1 U28644 ( .ip1(\LUT[86][0] ), .ip2(n27358), .op(n24575) );
  nand2_1 U28645 ( .ip1(n24576), .ip2(n24575), .op(n24577) );
  not_ab_or_c_or_d U28646 ( .ip1(n27363), .ip2(\LUT[87][0] ), .ip3(n24578), 
        .ip4(n24577), .op(n24579) );
  nor2_1 U28647 ( .ip1(n24579), .ip2(n27142), .op(n24618) );
  inv_1 U28648 ( .ip(n24580), .op(n24581) );
  nor2_1 U28649 ( .ip1(n24582), .ip2(n24581), .op(n27326) );
  inv_1 U28650 ( .ip(n24583), .op(n24585) );
  nor2_1 U28651 ( .ip1(n24585), .ip2(n24584), .op(n27317) );
  and2_1 U28652 ( .ip1(n27317), .ip2(\LUT[105][0] ), .op(n24603) );
  inv_1 U28653 ( .ip(n24586), .op(n24588) );
  nor2_1 U28654 ( .ip1(n24588), .ip2(n24587), .op(n27318) );
  nand2_1 U28655 ( .ip1(n27318), .ip2(\LUT[107][0] ), .op(n24601) );
  inv_1 U28656 ( .ip(n24589), .op(n24591) );
  nor2_1 U28657 ( .ip1(n24591), .ip2(n24590), .op(n27319) );
  nand2_1 U28658 ( .ip1(n27319), .ip2(\LUT[104][0] ), .op(n24600) );
  inv_1 U28659 ( .ip(n24592), .op(n24593) );
  nor2_1 U28660 ( .ip1(n24594), .ip2(n24593), .op(n27325) );
  nand2_1 U28661 ( .ip1(n27325), .ip2(\LUT[110][0] ), .op(n24599) );
  inv_1 U28662 ( .ip(n24595), .op(n24597) );
  nor2_1 U28663 ( .ip1(n24597), .ip2(n24596), .op(n27309) );
  nand2_1 U28664 ( .ip1(n27309), .ip2(\LUT[109][0] ), .op(n24598) );
  nand4_1 U28665 ( .ip1(n24601), .ip2(n24600), .ip3(n24599), .ip4(n24598), 
        .op(n24602) );
  not_ab_or_c_or_d U28666 ( .ip1(\LUT[102][0] ), .ip2(n27326), .ip3(n24603), 
        .ip4(n24602), .op(n24616) );
  inv_1 U28667 ( .ip(n24604), .op(n24605) );
  nor2_1 U28668 ( .ip1(n24606), .ip2(n24605), .op(n27370) );
  nand2_1 U28669 ( .ip1(n27370), .ip2(\LUT[100][0] ), .op(n24615) );
  inv_1 U28670 ( .ip(n24607), .op(n24609) );
  nor2_1 U28671 ( .ip1(n24609), .ip2(n24608), .op(n27328) );
  nand2_1 U28672 ( .ip1(n27328), .ip2(\LUT[101][0] ), .op(n24614) );
  inv_1 U28673 ( .ip(n24610), .op(n24611) );
  nor2_1 U28674 ( .ip1(n24612), .ip2(n24611), .op(n27327) );
  nand2_1 U28675 ( .ip1(n27327), .ip2(\LUT[103][0] ), .op(n24613) );
  nand4_1 U28676 ( .ip1(n24616), .ip2(n24615), .ip3(n24614), .ip4(n24613), 
        .op(n24617) );
  not_ab_or_c_or_d U28677 ( .ip1(\LUT[99][0] ), .ip2(n27156), .ip3(n24618), 
        .ip4(n24617), .op(n24619) );
  nor2_1 U28678 ( .ip1(n24619), .ip2(n27371), .op(n24647) );
  inv_1 U28679 ( .ip(n24620), .op(n24622) );
  nor2_1 U28680 ( .ip1(n24622), .ip2(n24621), .op(n27297) );
  inv_1 U28681 ( .ip(n24623), .op(n24624) );
  nor2_1 U28682 ( .ip1(n24625), .ip2(n24624), .op(n27582) );
  nand2_1 U28683 ( .ip1(n27582), .ip2(\LUT[115][0] ), .op(n24632) );
  inv_1 U28684 ( .ip(n24626), .op(n24627) );
  nor2_1 U28685 ( .ip1(n24628), .ip2(n24627), .op(n27298) );
  nand2_1 U28686 ( .ip1(n27298), .ip2(\LUT[117][0] ), .op(n24631) );
  nand2_1 U28687 ( .ip1(n27299), .ip2(\LUT[118][0] ), .op(n24630) );
  nand2_1 U28688 ( .ip1(n27300), .ip2(\LUT[119][0] ), .op(n24629) );
  nand4_1 U28689 ( .ip1(n24632), .ip2(n24631), .ip3(n24630), .ip4(n24629), 
        .op(n24633) );
  or2_1 U28690 ( .ip1(n27297), .ip2(n24633), .op(n24635) );
  or2_1 U28691 ( .ip1(\LUT[116][0] ), .ip2(n24633), .op(n24634) );
  nand2_1 U28692 ( .ip1(n24635), .ip2(n24634), .op(n24645) );
  inv_1 U28693 ( .ip(n24636), .op(n24637) );
  nor2_1 U28694 ( .ip1(n24638), .ip2(n24637), .op(n27583) );
  nand2_1 U28695 ( .ip1(n27583), .ip2(\LUT[113][0] ), .op(n24644) );
  nor2_1 U28696 ( .ip1(n26151), .ip2(n27371), .op(n27172) );
  nand2_1 U28697 ( .ip1(n27172), .ip2(\LUT[111][0] ), .op(n24643) );
  inv_1 U28698 ( .ip(n24639), .op(n24641) );
  nor2_1 U28699 ( .ip1(n24641), .ip2(n24640), .op(n27305) );
  nand2_1 U28700 ( .ip1(n27305), .ip2(\LUT[114][0] ), .op(n24642) );
  nand4_1 U28701 ( .ip1(n24645), .ip2(n24644), .ip3(n24643), .ip4(n24642), 
        .op(n24646) );
  not_ab_or_c_or_d U28702 ( .ip1(n27581), .ip2(\LUT[106][0] ), .ip3(n24647), 
        .ip4(n24646), .op(n24965) );
  inv_1 U28703 ( .ip(n24648), .op(n24650) );
  nor2_1 U28704 ( .ip1(n24650), .ip2(n24649), .op(n27390) );
  inv_1 U28705 ( .ip(n24651), .op(n24653) );
  nor2_1 U28706 ( .ip1(n24653), .ip2(n24652), .op(n27397) );
  inv_1 U28707 ( .ip(n24654), .op(n24655) );
  nor2_1 U28708 ( .ip1(n24656), .ip2(n24655), .op(n27542) );
  inv_1 U28709 ( .ip(n24657), .op(n24659) );
  nor2_1 U28710 ( .ip1(n24659), .ip2(n24658), .op(n27534) );
  and2_1 U28711 ( .ip1(n27534), .ip2(\LUT[65][0] ), .op(n24671) );
  inv_1 U28712 ( .ip(n24660), .op(n24662) );
  nor2_1 U28713 ( .ip1(n24662), .ip2(n24661), .op(n27548) );
  nand2_1 U28714 ( .ip1(n27548), .ip2(\LUT[67][0] ), .op(n24669) );
  nand2_1 U28715 ( .ip1(n27535), .ip2(\LUT[69][0] ), .op(n24668) );
  nand2_1 U28716 ( .ip1(n27536), .ip2(\LUT[70][0] ), .op(n24667) );
  inv_1 U28717 ( .ip(n24663), .op(n24664) );
  nor2_1 U28718 ( .ip1(n24665), .ip2(n24664), .op(n27537) );
  nand2_1 U28719 ( .ip1(n27537), .ip2(\LUT[68][0] ), .op(n24666) );
  nand4_1 U28720 ( .ip1(n24669), .ip2(n24668), .ip3(n24667), .ip4(n24666), 
        .op(n24670) );
  not_ab_or_c_or_d U28721 ( .ip1(n27542), .ip2(\LUT[66][0] ), .ip3(n24671), 
        .ip4(n24670), .op(n24682) );
  inv_1 U28722 ( .ip(n24672), .op(n24673) );
  nor2_1 U28723 ( .ip1(n24674), .ip2(n24673), .op(n27547) );
  nand2_1 U28724 ( .ip1(n27547), .ip2(\LUT[64][0] ), .op(n24681) );
  inv_1 U28725 ( .ip(n24675), .op(n24676) );
  nor2_1 U28726 ( .ip1(n24677), .ip2(n24676), .op(n27546) );
  nand2_1 U28727 ( .ip1(n27546), .ip2(\LUT[59][0] ), .op(n24680) );
  nor2_1 U28728 ( .ip1(n24687), .ip2(n24678), .op(n27556) );
  nand2_1 U28729 ( .ip1(n27556), .ip2(\LUT[63][0] ), .op(n24679) );
  nand4_1 U28730 ( .ip1(n24682), .ip2(n24681), .ip3(n24680), .ip4(n24679), 
        .op(n24699) );
  inv_1 U28731 ( .ip(n24683), .op(n24685) );
  nor2_1 U28732 ( .ip1(n24685), .ip2(n24684), .op(n27553) );
  nand2_1 U28733 ( .ip1(n27553), .ip2(\LUT[57][0] ), .op(n24697) );
  nor2_1 U28734 ( .ip1(n24687), .ip2(n24686), .op(n27563) );
  nand2_1 U28735 ( .ip1(n27563), .ip2(\LUT[62][0] ), .op(n24696) );
  inv_1 U28736 ( .ip(n24688), .op(n24689) );
  nor2_1 U28737 ( .ip1(n24690), .ip2(n24689), .op(n27555) );
  nand2_1 U28738 ( .ip1(n27555), .ip2(\LUT[61][0] ), .op(n24695) );
  inv_1 U28739 ( .ip(n24691), .op(n24693) );
  nor2_1 U28740 ( .ip1(n24693), .ip2(n24692), .op(n27554) );
  nand2_1 U28741 ( .ip1(n27554), .ip2(\LUT[60][0] ), .op(n24694) );
  nand4_1 U28742 ( .ip1(n24697), .ip2(n24696), .ip3(n24695), .ip4(n24694), 
        .op(n24698) );
  not_ab_or_c_or_d U28743 ( .ip1(n27397), .ip2(\LUT[58][0] ), .ip3(n24699), 
        .ip4(n24698), .op(n24700) );
  inv_1 U28744 ( .ip(n27567), .op(n27265) );
  or2_1 U28745 ( .ip1(n24700), .ip2(n27265), .op(n24906) );
  inv_1 U28746 ( .ip(n24701), .op(n24702) );
  nor2_1 U28747 ( .ip1(n24703), .ip2(n24702), .op(n27459) );
  nand2_1 U28748 ( .ip1(\LUT[27][0] ), .ip2(n27398), .op(n24708) );
  nand2_1 U28749 ( .ip1(n27400), .ip2(\LUT[28][0] ), .op(n24707) );
  inv_1 U28750 ( .ip(n24704), .op(n24716) );
  nor2_1 U28751 ( .ip1(n24716), .ip2(n24705), .op(n27405) );
  nand2_1 U28752 ( .ip1(n27405), .ip2(\LUT[25][0] ), .op(n24706) );
  nand3_1 U28753 ( .ip1(n24708), .ip2(n24707), .ip3(n24706), .op(n24721) );
  inv_1 U28754 ( .ip(n24709), .op(n24711) );
  nor2_1 U28755 ( .ip1(n24711), .ip2(n24710), .op(n27404) );
  nand2_1 U28756 ( .ip1(\LUT[24][0] ), .ip2(n27404), .op(n24719) );
  inv_1 U28757 ( .ip(n24712), .op(n24713) );
  nor2_1 U28758 ( .ip1(n24714), .ip2(n24713), .op(n27406) );
  nand2_1 U28759 ( .ip1(n27406), .ip2(\LUT[23][0] ), .op(n24718) );
  nor2_1 U28760 ( .ip1(n24716), .ip2(n24715), .op(n27399) );
  nand2_1 U28761 ( .ip1(n27399), .ip2(\LUT[26][0] ), .op(n24717) );
  nand3_1 U28762 ( .ip1(n24719), .ip2(n24718), .ip3(n24717), .op(n24720) );
  not_ab_or_c_or_d U28763 ( .ip1(n27459), .ip2(\LUT[17][0] ), .ip3(n24721), 
        .ip4(n24720), .op(n24799) );
  inv_1 U28764 ( .ip(n24722), .op(n24723) );
  nor2_1 U28765 ( .ip1(n24724), .ip2(n24723), .op(n27458) );
  inv_1 U28766 ( .ip(n24725), .op(n24728) );
  nor2_1 U28767 ( .ip1(n24728), .ip2(n24726), .op(n27413) );
  nand2_1 U28768 ( .ip1(\LUT[2][0] ), .ip2(n27413), .op(n24730) );
  nor2_1 U28769 ( .ip1(n24728), .ip2(n24727), .op(n27414) );
  nand2_1 U28770 ( .ip1(\LUT[3][0] ), .ip2(n27414), .op(n24729) );
  nand2_1 U28771 ( .ip1(n24730), .ip2(n24729), .op(n24771) );
  inv_1 U28772 ( .ip(n24731), .op(n24732) );
  nor2_1 U28773 ( .ip1(n24733), .ip2(n24732), .op(n27418) );
  inv_1 U28774 ( .ip(n24734), .op(n24751) );
  nor2_1 U28775 ( .ip1(n24751), .ip2(n24735), .op(n27417) );
  nand2_1 U28776 ( .ip1(n27417), .ip2(\LUT[7][0] ), .op(n24741) );
  inv_1 U28777 ( .ip(n24736), .op(n24749) );
  nor2_1 U28778 ( .ip1(n24749), .ip2(n24737), .op(n27427) );
  nand2_1 U28779 ( .ip1(n27427), .ip2(\LUT[12][0] ), .op(n24740) );
  nand2_1 U28780 ( .ip1(n27419), .ip2(\LUT[14][0] ), .op(n24739) );
  nand2_1 U28781 ( .ip1(n27420), .ip2(\LUT[13][0] ), .op(n24738) );
  nand4_1 U28782 ( .ip1(n24741), .ip2(n24740), .ip3(n24739), .ip4(n24738), 
        .op(n24757) );
  inv_1 U28783 ( .ip(n24742), .op(n24744) );
  nor2_1 U28784 ( .ip1(n24744), .ip2(n24743), .op(n27426) );
  nand2_1 U28785 ( .ip1(n27426), .ip2(\LUT[8][0] ), .op(n24755) );
  inv_1 U28786 ( .ip(n24745), .op(n24747) );
  nor2_1 U28787 ( .ip1(n24747), .ip2(n24746), .op(n27425) );
  nand2_1 U28788 ( .ip1(n27425), .ip2(\LUT[10][0] ), .op(n24754) );
  nor2_1 U28789 ( .ip1(n24749), .ip2(n24748), .op(n27435) );
  nand2_1 U28790 ( .ip1(n27435), .ip2(\LUT[11][0] ), .op(n24753) );
  nor2_1 U28791 ( .ip1(n24751), .ip2(n24750), .op(n27428) );
  nand2_1 U28792 ( .ip1(n27428), .ip2(\LUT[6][0] ), .op(n24752) );
  nand4_1 U28793 ( .ip1(n24755), .ip2(n24754), .ip3(n24753), .ip4(n24752), 
        .op(n24756) );
  not_ab_or_c_or_d U28794 ( .ip1(n27418), .ip2(\LUT[9][0] ), .ip3(n24757), 
        .ip4(n24756), .op(n24769) );
  inv_1 U28795 ( .ip(n24758), .op(n24759) );
  nor2_1 U28796 ( .ip1(n24760), .ip2(n24759), .op(n27445) );
  nand2_1 U28797 ( .ip1(n27445), .ip2(\LUT[1][0] ), .op(n24768) );
  inv_1 U28798 ( .ip(n24761), .op(n24762) );
  nor2_1 U28799 ( .ip1(n24765), .ip2(n24762), .op(n27438) );
  nand2_1 U28800 ( .ip1(n27438), .ip2(\LUT[5][0] ), .op(n24767) );
  inv_1 U28801 ( .ip(n24763), .op(n24764) );
  nor2_1 U28802 ( .ip1(n24765), .ip2(n24764), .op(n27437) );
  nand2_1 U28803 ( .ip1(n27437), .ip2(\LUT[4][0] ), .op(n24766) );
  nand4_1 U28804 ( .ip1(n24769), .ip2(n24768), .ip3(n24767), .ip4(n24766), 
        .op(n24770) );
  not_ab_or_c_or_d U28805 ( .ip1(n27436), .ip2(\LUT[0][0] ), .ip3(n24771), 
        .ip4(n24770), .op(n24773) );
  inv_1 U28806 ( .ip(n24772), .op(n27446) );
  nor2_1 U28807 ( .ip1(n24773), .ip2(n27446), .op(n24789) );
  inv_1 U28808 ( .ip(n24774), .op(n24775) );
  nor2_1 U28809 ( .ip1(n24776), .ip2(n24775), .op(n27448) );
  nand2_1 U28810 ( .ip1(n27448), .ip2(\LUT[18][0] ), .op(n24787) );
  inv_1 U28811 ( .ip(n24777), .op(n24780) );
  nor2_1 U28812 ( .ip1(n24780), .ip2(n24778), .op(n27450) );
  nand2_1 U28813 ( .ip1(n27450), .ip2(\LUT[21][0] ), .op(n24786) );
  nor2_1 U28814 ( .ip1(n24780), .ip2(n24779), .op(n27449) );
  nand2_1 U28815 ( .ip1(n27449), .ip2(\LUT[20][0] ), .op(n24785) );
  inv_1 U28816 ( .ip(n24781), .op(n24783) );
  nor2_1 U28817 ( .ip1(n24783), .ip2(n24782), .op(n27451) );
  nand2_1 U28818 ( .ip1(n27451), .ip2(\LUT[16][0] ), .op(n24784) );
  nand4_1 U28819 ( .ip1(n24787), .ip2(n24786), .ip3(n24785), .ip4(n24784), 
        .op(n24788) );
  not_ab_or_c_or_d U28820 ( .ip1(\LUT[15][0] ), .ip2(n27458), .ip3(n24789), 
        .ip4(n24788), .op(n24798) );
  inv_1 U28821 ( .ip(n24790), .op(n24792) );
  nor2_1 U28822 ( .ip1(n24792), .ip2(n24791), .op(n27460) );
  nand2_1 U28823 ( .ip1(n27460), .ip2(\LUT[19][0] ), .op(n24797) );
  inv_1 U28824 ( .ip(n24793), .op(n24795) );
  nor2_1 U28825 ( .ip1(n24795), .ip2(n24794), .op(n27412) );
  nand2_1 U28826 ( .ip1(n27412), .ip2(\LUT[22][0] ), .op(n24796) );
  nand4_1 U28827 ( .ip1(n24799), .ip2(n24798), .ip3(n24797), .ip4(n24796), 
        .op(n24903) );
  inv_1 U28828 ( .ip(n24800), .op(n24801) );
  nor2_1 U28829 ( .ip1(n24802), .ip2(n24801), .op(n27527) );
  and2_1 U28830 ( .ip1(n24840), .ip2(n24803), .op(n27499) );
  nand2_1 U28831 ( .ip1(n27499), .ip2(\LUT[49][0] ), .op(n24815) );
  inv_1 U28832 ( .ip(n24804), .op(n24805) );
  nor2_1 U28833 ( .ip1(n24806), .ip2(n24805), .op(n27498) );
  nand2_1 U28834 ( .ip1(n27498), .ip2(\LUT[48][0] ), .op(n24814) );
  inv_1 U28835 ( .ip(n24807), .op(n24808) );
  nor2_1 U28836 ( .ip1(n24809), .ip2(n24808), .op(n27501) );
  nand2_1 U28837 ( .ip1(n27501), .ip2(\LUT[52][0] ), .op(n24813) );
  inv_1 U28838 ( .ip(n24810), .op(n24811) );
  nor2_1 U28839 ( .ip1(n24826), .ip2(n24811), .op(n27507) );
  nand2_1 U28840 ( .ip1(n27507), .ip2(\LUT[54][0] ), .op(n24812) );
  nand4_1 U28841 ( .ip1(n24815), .ip2(n24814), .ip3(n24813), .ip4(n24812), 
        .op(n24848) );
  inv_1 U28842 ( .ip(n24816), .op(n24818) );
  nor2_1 U28843 ( .ip1(n24818), .ip2(n24817), .op(n27520) );
  inv_1 U28844 ( .ip(n24819), .op(n24839) );
  nor2_1 U28845 ( .ip1(n24839), .ip2(n24820), .op(n27518) );
  and2_1 U28846 ( .ip1(n27518), .ip2(\LUT[44][0] ), .op(n24834) );
  inv_1 U28847 ( .ip(n24821), .op(n24823) );
  nor2_1 U28848 ( .ip1(n24823), .ip2(n24822), .op(n27510) );
  nand2_1 U28849 ( .ip1(n27510), .ip2(\LUT[51][0] ), .op(n24832) );
  inv_1 U28850 ( .ip(n24824), .op(n24825) );
  nor2_1 U28851 ( .ip1(n24826), .ip2(n24825), .op(n27500) );
  nand2_1 U28852 ( .ip1(n27500), .ip2(\LUT[53][0] ), .op(n24831) );
  inv_1 U28853 ( .ip(n24827), .op(n27508) );
  nand2_1 U28854 ( .ip1(n27508), .ip2(\LUT[55][0] ), .op(n24830) );
  inv_1 U28855 ( .ip(n24828), .op(n27509) );
  nand2_1 U28856 ( .ip1(n27509), .ip2(\LUT[56][0] ), .op(n24829) );
  nand4_1 U28857 ( .ip1(n24832), .ip2(n24831), .ip3(n24830), .ip4(n24829), 
        .op(n24833) );
  not_ab_or_c_or_d U28858 ( .ip1(\LUT[47][0] ), .ip2(n27520), .ip3(n24834), 
        .ip4(n24833), .op(n24846) );
  inv_1 U28859 ( .ip(n24835), .op(n24836) );
  nor2_1 U28860 ( .ip1(n24837), .ip2(n24836), .op(n27519) );
  nand2_1 U28861 ( .ip1(n27519), .ip2(\LUT[43][0] ), .op(n24845) );
  nor2_1 U28862 ( .ip1(n24839), .ip2(n24838), .op(n27506) );
  nand2_1 U28863 ( .ip1(n27506), .ip2(\LUT[45][0] ), .op(n24844) );
  inv_1 U28864 ( .ip(n24840), .op(n24841) );
  nor2_1 U28865 ( .ip1(n24842), .ip2(n24841), .op(n27517) );
  nand2_1 U28866 ( .ip1(n27517), .ip2(\LUT[50][0] ), .op(n24843) );
  nand4_1 U28867 ( .ip1(n24846), .ip2(n24845), .ip3(n24844), .ip4(n24843), 
        .op(n24847) );
  not_ab_or_c_or_d U28868 ( .ip1(n27527), .ip2(\LUT[46][0] ), .ip3(n24848), 
        .ip4(n24847), .op(n24849) );
  inv_1 U28869 ( .ip(n26760), .op(n27528) );
  nor2_1 U28870 ( .ip1(n24849), .ip2(n27528), .op(n24902) );
  inv_1 U28871 ( .ip(n24850), .op(n24851) );
  nor2_1 U28872 ( .ip1(n24852), .ip2(n24851), .op(n27495) );
  inv_1 U28873 ( .ip(n24853), .op(n24856) );
  nor2_1 U28874 ( .ip1(n24856), .ip2(n24854), .op(n27465) );
  nand2_1 U28875 ( .ip1(\LUT[31][0] ), .ip2(n27465), .op(n24858) );
  nor2_1 U28876 ( .ip1(n24856), .ip2(n24855), .op(n27466) );
  nand2_1 U28877 ( .ip1(\LUT[30][0] ), .ip2(n27466), .op(n24857) );
  nand2_1 U28878 ( .ip1(n24858), .ip2(n24857), .op(n24899) );
  inv_1 U28879 ( .ip(n24859), .op(n24861) );
  nor2_1 U28880 ( .ip1(n24861), .ip2(n24860), .op(n27485) );
  inv_1 U28881 ( .ip(n24862), .op(n24864) );
  nor2_1 U28882 ( .ip1(n24864), .ip2(n24863), .op(n27470) );
  nand2_1 U28883 ( .ip1(n27470), .ip2(\LUT[38][0] ), .op(n24873) );
  inv_1 U28884 ( .ip(n24865), .op(n24866) );
  nor2_1 U28885 ( .ip1(n24867), .ip2(n24866), .op(n27469) );
  nand2_1 U28886 ( .ip1(n27469), .ip2(\LUT[39][0] ), .op(n24872) );
  inv_1 U28887 ( .ip(n24868), .op(n27471) );
  nand2_1 U28888 ( .ip1(n27471), .ip2(\LUT[41][0] ), .op(n24871) );
  inv_1 U28889 ( .ip(n24869), .op(n27472) );
  nand2_1 U28890 ( .ip1(n27472), .ip2(\LUT[42][0] ), .op(n24870) );
  nand4_1 U28891 ( .ip1(n24873), .ip2(n24872), .ip3(n24871), .ip4(n24870), 
        .op(n24886) );
  inv_1 U28892 ( .ip(n24874), .op(n24876) );
  nor2_1 U28893 ( .ip1(n24876), .ip2(n24875), .op(n27477) );
  nand2_1 U28894 ( .ip1(\LUT[36][0] ), .ip2(n27477), .op(n24884) );
  inv_1 U28895 ( .ip(n24877), .op(n24879) );
  nor2_1 U28896 ( .ip1(n24879), .ip2(n24878), .op(n27478) );
  nand2_1 U28897 ( .ip1(n27478), .ip2(\LUT[37][0] ), .op(n24883) );
  inv_1 U28898 ( .ip(n24880), .op(n24881) );
  nor2_1 U28899 ( .ip1(n24891), .ip2(n24881), .op(n27479) );
  nand2_1 U28900 ( .ip1(n27479), .ip2(\LUT[32][0] ), .op(n24882) );
  nand3_1 U28901 ( .ip1(n24884), .ip2(n24883), .ip3(n24882), .op(n24885) );
  not_ab_or_c_or_d U28902 ( .ip1(n27485), .ip2(\LUT[40][0] ), .ip3(n24886), 
        .ip4(n24885), .op(n24897) );
  inv_1 U28903 ( .ip(n24887), .op(n24893) );
  nor2_1 U28904 ( .ip1(n24893), .ip2(n24888), .op(n27486) );
  nand2_1 U28905 ( .ip1(n27486), .ip2(\LUT[34][0] ), .op(n24896) );
  inv_1 U28906 ( .ip(n24889), .op(n24890) );
  nor2_1 U28907 ( .ip1(n24891), .ip2(n24890), .op(n27488) );
  nand2_1 U28908 ( .ip1(n27488), .ip2(\LUT[33][0] ), .op(n24895) );
  nor2_1 U28909 ( .ip1(n24893), .ip2(n24892), .op(n27487) );
  nand2_1 U28910 ( .ip1(n27487), .ip2(\LUT[35][0] ), .op(n24894) );
  nand4_1 U28911 ( .ip1(n24897), .ip2(n24896), .ip3(n24895), .ip4(n24894), 
        .op(n24898) );
  not_ab_or_c_or_d U28912 ( .ip1(n27495), .ip2(\LUT[29][0] ), .ip3(n24899), 
        .ip4(n24898), .op(n24900) );
  nor2_1 U28913 ( .ip1(n24900), .ip2(n27496), .op(n24901) );
  not_ab_or_c_or_d U28914 ( .ip1(n27533), .ip2(n24903), .ip3(n24902), .ip4(
        n24901), .op(n24904) );
  or2_1 U28915 ( .ip1(n24904), .ip2(n27265), .op(n24905) );
  nand2_1 U28916 ( .ip1(n24906), .ip2(n24905), .op(n24946) );
  inv_1 U28917 ( .ip(n24907), .op(n24908) );
  nor2_1 U28918 ( .ip1(n24909), .ip2(n24908), .op(n27391) );
  nand2_1 U28919 ( .ip1(n27391), .ip2(\LUT[75][0] ), .op(n24944) );
  inv_1 U28920 ( .ip(n24910), .op(n24911) );
  nor2_1 U28921 ( .ip1(n24912), .ip2(n24911), .op(n27389) );
  inv_1 U28922 ( .ip(n24913), .op(n24914) );
  nor2_1 U28923 ( .ip1(n24915), .ip2(n24914), .op(n27373) );
  nand2_1 U28924 ( .ip1(n27373), .ip2(\LUT[82][0] ), .op(n24924) );
  inv_1 U28925 ( .ip(n24916), .op(n24918) );
  nor2_1 U28926 ( .ip1(n24918), .ip2(n24917), .op(n27374) );
  nand2_1 U28927 ( .ip1(n27374), .ip2(\LUT[81][0] ), .op(n24923) );
  inv_1 U28928 ( .ip(n24919), .op(n27376) );
  nand2_1 U28929 ( .ip1(n27376), .ip2(\LUT[83][0] ), .op(n24922) );
  inv_1 U28930 ( .ip(n24920), .op(n27375) );
  nand2_1 U28931 ( .ip1(n27375), .ip2(\LUT[84][0] ), .op(n24921) );
  nand4_1 U28932 ( .ip1(n24924), .ip2(n24923), .ip3(n24922), .ip4(n24921), 
        .op(n24938) );
  inv_1 U28933 ( .ip(n24925), .op(n24926) );
  nor2_1 U28934 ( .ip1(n24927), .ip2(n24926), .op(n27381) );
  nand2_1 U28935 ( .ip1(n27381), .ip2(\LUT[78][0] ), .op(n24936) );
  inv_1 U28936 ( .ip(n24928), .op(n24930) );
  nor2_1 U28937 ( .ip1(n24930), .ip2(n24929), .op(n27382) );
  nand2_1 U28938 ( .ip1(n27382), .ip2(\LUT[79][0] ), .op(n24935) );
  inv_1 U28939 ( .ip(n24931), .op(n24932) );
  nor2_1 U28940 ( .ip1(n24933), .ip2(n24932), .op(n27383) );
  nand2_1 U28941 ( .ip1(n27383), .ip2(\LUT[77][0] ), .op(n24934) );
  nand3_1 U28942 ( .ip1(n24936), .ip2(n24935), .ip3(n24934), .op(n24937) );
  not_ab_or_c_or_d U28943 ( .ip1(n27389), .ip2(\LUT[80][0] ), .ip3(n24938), 
        .ip4(n24937), .op(n24943) );
  inv_1 U28944 ( .ip(n24939), .op(n24941) );
  nor2_1 U28945 ( .ip1(n24941), .ip2(n24940), .op(n27392) );
  nand2_1 U28946 ( .ip1(n27392), .ip2(\LUT[74][0] ), .op(n24942) );
  nand3_1 U28947 ( .ip1(n24944), .ip2(n24943), .ip3(n24942), .op(n24945) );
  not_ab_or_c_or_d U28948 ( .ip1(n27390), .ip2(\LUT[76][0] ), .ip3(n24946), 
        .ip4(n24945), .op(n24957) );
  inv_1 U28949 ( .ip(n24947), .op(n24948) );
  nor2_1 U28950 ( .ip1(n24949), .ip2(n24948), .op(n27576) );
  nand2_1 U28951 ( .ip1(n27576), .ip2(\LUT[71][0] ), .op(n24956) );
  inv_1 U28952 ( .ip(n24950), .op(n24953) );
  nor2_1 U28953 ( .ip1(n24953), .ip2(n24951), .op(n27570) );
  nand2_1 U28954 ( .ip1(n27570), .ip2(\LUT[72][0] ), .op(n24955) );
  nor2_1 U28955 ( .ip1(n24953), .ip2(n24952), .op(n27569) );
  nand2_1 U28956 ( .ip1(n27569), .ip2(\LUT[73][0] ), .op(n24954) );
  nand4_1 U28957 ( .ip1(n24957), .ip2(n24956), .ip3(n24955), .ip4(n24954), 
        .op(n24958) );
  nand2_1 U28958 ( .ip1(n27288), .ip2(n24958), .op(n24964) );
  nor2_1 U28959 ( .ip1(n26152), .ip2(n27371), .op(n27289) );
  nand2_1 U28960 ( .ip1(n27289), .ip2(\LUT[112][0] ), .op(n24963) );
  inv_1 U28961 ( .ip(n24959), .op(n24961) );
  nand2_1 U28962 ( .ip1(n24961), .ip2(n24960), .op(n26155) );
  nor2_1 U28963 ( .ip1(n27371), .ip2(n26155), .op(n27165) );
  nand2_1 U28964 ( .ip1(n27165), .ip2(\LUT[108][0] ), .op(n24962) );
  nand4_1 U28965 ( .ip1(n24965), .ip2(n24964), .ip3(n24963), .ip4(n24962), 
        .op(n24966) );
  nand2_1 U28966 ( .ip1(n27589), .ip2(n24966), .op(n24972) );
  or2_1 U28967 ( .ip1(done), .ip2(reset), .op(n24969) );
  or2_1 U28968 ( .ip1(n24967), .ip2(reset), .op(n24968) );
  nand2_1 U28969 ( .ip1(n24969), .ip2(n24968), .op(n24970) );
  or2_1 U28970 ( .ip1(we), .ip2(n24970), .op(n27590) );
  nand2_1 U28971 ( .ip1(sig_out[0]), .ip2(n27590), .op(n24971) );
  nand2_1 U28972 ( .ip1(n24972), .ip2(n24971), .op(n13465) );
  nand2_1 U28973 ( .ip1(n27333), .ip2(\LUT[95][1] ), .op(n24976) );
  nand2_1 U28974 ( .ip1(n27334), .ip2(\LUT[94][1] ), .op(n24975) );
  nand2_1 U28975 ( .ip1(n27336), .ip2(\LUT[97][1] ), .op(n24974) );
  nand2_1 U28976 ( .ip1(n27335), .ip2(\LUT[98][1] ), .op(n24973) );
  nand4_1 U28977 ( .ip1(n24976), .ip2(n24975), .ip3(n24974), .ip4(n24973), 
        .op(n24981) );
  nand2_1 U28978 ( .ip1(n27341), .ip2(\LUT[93][1] ), .op(n24979) );
  nand2_1 U28979 ( .ip1(n27342), .ip2(\LUT[92][1] ), .op(n24978) );
  nand2_1 U28980 ( .ip1(n27343), .ip2(\LUT[91][1] ), .op(n24977) );
  nand3_1 U28981 ( .ip1(n24979), .ip2(n24978), .ip3(n24977), .op(n24980) );
  not_ab_or_c_or_d U28982 ( .ip1(n27349), .ip2(\LUT[96][1] ), .ip3(n24981), 
        .ip4(n24980), .op(n24985) );
  nand2_1 U28983 ( .ip1(n27350), .ip2(\LUT[89][1] ), .op(n24984) );
  nand2_1 U28984 ( .ip1(n27351), .ip2(\LUT[90][1] ), .op(n24983) );
  nand2_1 U28985 ( .ip1(n27352), .ip2(\LUT[88][1] ), .op(n24982) );
  nand4_1 U28986 ( .ip1(n24985), .ip2(n24984), .ip3(n24983), .ip4(n24982), 
        .op(n24989) );
  nand2_1 U28987 ( .ip1(\LUT[85][1] ), .ip2(n27357), .op(n24987) );
  nand2_1 U28988 ( .ip1(\LUT[86][1] ), .ip2(n27358), .op(n24986) );
  nand2_1 U28989 ( .ip1(n24987), .ip2(n24986), .op(n24988) );
  not_ab_or_c_or_d U28990 ( .ip1(n27363), .ip2(\LUT[87][1] ), .ip3(n24989), 
        .ip4(n24988), .op(n24990) );
  nor2_1 U28991 ( .ip1(n24990), .ip2(n27142), .op(n25002) );
  and2_1 U28992 ( .ip1(n27317), .ip2(\LUT[105][1] ), .op(n24996) );
  nand2_1 U28993 ( .ip1(n27318), .ip2(\LUT[107][1] ), .op(n24994) );
  nand2_1 U28994 ( .ip1(n27319), .ip2(\LUT[104][1] ), .op(n24993) );
  nand2_1 U28995 ( .ip1(n27309), .ip2(\LUT[109][1] ), .op(n24992) );
  nand2_1 U28996 ( .ip1(n27325), .ip2(\LUT[110][1] ), .op(n24991) );
  nand4_1 U28997 ( .ip1(n24994), .ip2(n24993), .ip3(n24992), .ip4(n24991), 
        .op(n24995) );
  not_ab_or_c_or_d U28998 ( .ip1(\LUT[102][1] ), .ip2(n27326), .ip3(n24996), 
        .ip4(n24995), .op(n25000) );
  nand2_1 U28999 ( .ip1(n27370), .ip2(\LUT[100][1] ), .op(n24999) );
  nand2_1 U29000 ( .ip1(n27328), .ip2(\LUT[101][1] ), .op(n24998) );
  nand2_1 U29001 ( .ip1(n27327), .ip2(\LUT[103][1] ), .op(n24997) );
  nand4_1 U29002 ( .ip1(n25000), .ip2(n24999), .ip3(n24998), .ip4(n24997), 
        .op(n25001) );
  not_ab_or_c_or_d U29003 ( .ip1(\LUT[99][1] ), .ip2(n27156), .ip3(n25002), 
        .ip4(n25001), .op(n25003) );
  nor2_1 U29004 ( .ip1(n25003), .ip2(n27371), .op(n25016) );
  nand2_1 U29005 ( .ip1(n27305), .ip2(\LUT[114][1] ), .op(n25007) );
  nand2_1 U29006 ( .ip1(n27298), .ip2(\LUT[117][1] ), .op(n25006) );
  nand2_1 U29007 ( .ip1(n27299), .ip2(\LUT[118][1] ), .op(n25005) );
  nand2_1 U29008 ( .ip1(n27300), .ip2(\LUT[119][1] ), .op(n25004) );
  nand4_1 U29009 ( .ip1(n25007), .ip2(n25006), .ip3(n25005), .ip4(n25004), 
        .op(n25008) );
  or2_1 U29010 ( .ip1(n27297), .ip2(n25008), .op(n25010) );
  or2_1 U29011 ( .ip1(\LUT[116][1] ), .ip2(n25008), .op(n25009) );
  nand2_1 U29012 ( .ip1(n25010), .ip2(n25009), .op(n25014) );
  nand2_1 U29013 ( .ip1(n27289), .ip2(\LUT[112][1] ), .op(n25013) );
  nand2_1 U29014 ( .ip1(n27583), .ip2(\LUT[113][1] ), .op(n25012) );
  nand2_1 U29015 ( .ip1(n27582), .ip2(\LUT[115][1] ), .op(n25011) );
  nand4_1 U29016 ( .ip1(n25014), .ip2(n25013), .ip3(n25012), .ip4(n25011), 
        .op(n25015) );
  not_ab_or_c_or_d U29017 ( .ip1(n27581), .ip2(\LUT[106][1] ), .ip3(n25016), 
        .ip4(n25015), .op(n25134) );
  and2_1 U29018 ( .ip1(n27548), .ip2(\LUT[67][1] ), .op(n25022) );
  nand2_1 U29019 ( .ip1(n27534), .ip2(\LUT[65][1] ), .op(n25020) );
  nand2_1 U29020 ( .ip1(n27535), .ip2(\LUT[69][1] ), .op(n25019) );
  nand2_1 U29021 ( .ip1(n27536), .ip2(\LUT[70][1] ), .op(n25018) );
  nand2_1 U29022 ( .ip1(n27537), .ip2(\LUT[68][1] ), .op(n25017) );
  nand4_1 U29023 ( .ip1(n25020), .ip2(n25019), .ip3(n25018), .ip4(n25017), 
        .op(n25021) );
  not_ab_or_c_or_d U29024 ( .ip1(n27542), .ip2(\LUT[66][1] ), .ip3(n25022), 
        .ip4(n25021), .op(n25026) );
  nand2_1 U29025 ( .ip1(n27546), .ip2(\LUT[59][1] ), .op(n25025) );
  nand2_1 U29026 ( .ip1(n27563), .ip2(\LUT[62][1] ), .op(n25024) );
  nand2_1 U29027 ( .ip1(n27547), .ip2(\LUT[64][1] ), .op(n25023) );
  nand4_1 U29028 ( .ip1(n25026), .ip2(n25025), .ip3(n25024), .ip4(n25023), 
        .op(n25032) );
  nand2_1 U29029 ( .ip1(n27397), .ip2(\LUT[58][1] ), .op(n25030) );
  nand2_1 U29030 ( .ip1(n27556), .ip2(\LUT[63][1] ), .op(n25029) );
  nand2_1 U29031 ( .ip1(n27555), .ip2(\LUT[61][1] ), .op(n25028) );
  nand2_1 U29032 ( .ip1(n27554), .ip2(\LUT[60][1] ), .op(n25027) );
  nand4_1 U29033 ( .ip1(n25030), .ip2(n25029), .ip3(n25028), .ip4(n25027), 
        .op(n25031) );
  not_ab_or_c_or_d U29034 ( .ip1(n27553), .ip2(\LUT[57][1] ), .ip3(n25032), 
        .ip4(n25031), .op(n25033) );
  or2_1 U29035 ( .ip1(n25033), .ip2(n27265), .op(n25111) );
  nand2_1 U29036 ( .ip1(\LUT[27][1] ), .ip2(n27398), .op(n25036) );
  nand2_1 U29037 ( .ip1(n27400), .ip2(\LUT[28][1] ), .op(n25035) );
  nand2_1 U29038 ( .ip1(n27399), .ip2(\LUT[26][1] ), .op(n25034) );
  nand3_1 U29039 ( .ip1(n25036), .ip2(n25035), .ip3(n25034), .op(n25041) );
  nand2_1 U29040 ( .ip1(\LUT[24][1] ), .ip2(n27404), .op(n25039) );
  nand2_1 U29041 ( .ip1(n27405), .ip2(\LUT[25][1] ), .op(n25038) );
  nand2_1 U29042 ( .ip1(n27406), .ip2(\LUT[23][1] ), .op(n25037) );
  nand3_1 U29043 ( .ip1(n25039), .ip2(n25038), .ip3(n25037), .op(n25040) );
  not_ab_or_c_or_d U29044 ( .ip1(n27412), .ip2(\LUT[22][1] ), .ip3(n25041), 
        .ip4(n25040), .op(n25070) );
  nand2_1 U29045 ( .ip1(\LUT[2][1] ), .ip2(n27413), .op(n25043) );
  nand2_1 U29046 ( .ip1(\LUT[3][1] ), .ip2(n27414), .op(n25042) );
  nand2_1 U29047 ( .ip1(n25043), .ip2(n25042), .op(n25059) );
  nand2_1 U29048 ( .ip1(n27418), .ip2(\LUT[9][1] ), .op(n25047) );
  nand2_1 U29049 ( .ip1(n27417), .ip2(\LUT[7][1] ), .op(n25046) );
  nand2_1 U29050 ( .ip1(n27420), .ip2(\LUT[13][1] ), .op(n25045) );
  nand2_1 U29051 ( .ip1(n27419), .ip2(\LUT[14][1] ), .op(n25044) );
  nand4_1 U29052 ( .ip1(n25047), .ip2(n25046), .ip3(n25045), .ip4(n25044), 
        .op(n25053) );
  nand2_1 U29053 ( .ip1(n27426), .ip2(\LUT[8][1] ), .op(n25051) );
  nand2_1 U29054 ( .ip1(n27425), .ip2(\LUT[10][1] ), .op(n25050) );
  nand2_1 U29055 ( .ip1(n27427), .ip2(\LUT[12][1] ), .op(n25049) );
  nand2_1 U29056 ( .ip1(n27428), .ip2(\LUT[6][1] ), .op(n25048) );
  nand4_1 U29057 ( .ip1(n25051), .ip2(n25050), .ip3(n25049), .ip4(n25048), 
        .op(n25052) );
  not_ab_or_c_or_d U29058 ( .ip1(n27435), .ip2(\LUT[11][1] ), .ip3(n25053), 
        .ip4(n25052), .op(n25057) );
  nand2_1 U29059 ( .ip1(n27445), .ip2(\LUT[1][1] ), .op(n25056) );
  nand2_1 U29060 ( .ip1(n27438), .ip2(\LUT[5][1] ), .op(n25055) );
  nand2_1 U29061 ( .ip1(n27437), .ip2(\LUT[4][1] ), .op(n25054) );
  nand4_1 U29062 ( .ip1(n25057), .ip2(n25056), .ip3(n25055), .ip4(n25054), 
        .op(n25058) );
  not_ab_or_c_or_d U29063 ( .ip1(n27436), .ip2(\LUT[0][1] ), .ip3(n25059), 
        .ip4(n25058), .op(n25060) );
  nor2_1 U29064 ( .ip1(n25060), .ip2(n27446), .op(n25066) );
  nand2_1 U29065 ( .ip1(n27448), .ip2(\LUT[18][1] ), .op(n25064) );
  nand2_1 U29066 ( .ip1(n27450), .ip2(\LUT[21][1] ), .op(n25063) );
  nand2_1 U29067 ( .ip1(n27449), .ip2(\LUT[20][1] ), .op(n25062) );
  nand2_1 U29068 ( .ip1(n27451), .ip2(\LUT[16][1] ), .op(n25061) );
  nand4_1 U29069 ( .ip1(n25064), .ip2(n25063), .ip3(n25062), .ip4(n25061), 
        .op(n25065) );
  not_ab_or_c_or_d U29070 ( .ip1(\LUT[15][1] ), .ip2(n27458), .ip3(n25066), 
        .ip4(n25065), .op(n25069) );
  nand2_1 U29071 ( .ip1(n27459), .ip2(\LUT[17][1] ), .op(n25068) );
  nand2_1 U29072 ( .ip1(n27460), .ip2(\LUT[19][1] ), .op(n25067) );
  nand4_1 U29073 ( .ip1(n25070), .ip2(n25069), .ip3(n25068), .ip4(n25067), 
        .op(n25108) );
  nand2_1 U29074 ( .ip1(\LUT[31][1] ), .ip2(n27465), .op(n25072) );
  nand2_1 U29075 ( .ip1(\LUT[30][1] ), .ip2(n27466), .op(n25071) );
  nand2_1 U29076 ( .ip1(n25072), .ip2(n25071), .op(n25087) );
  nand2_1 U29077 ( .ip1(n27470), .ip2(\LUT[38][1] ), .op(n25076) );
  nand2_1 U29078 ( .ip1(n27469), .ip2(\LUT[39][1] ), .op(n25075) );
  nand2_1 U29079 ( .ip1(n27472), .ip2(\LUT[42][1] ), .op(n25074) );
  nand2_1 U29080 ( .ip1(n27471), .ip2(\LUT[41][1] ), .op(n25073) );
  nand4_1 U29081 ( .ip1(n25076), .ip2(n25075), .ip3(n25074), .ip4(n25073), 
        .op(n25081) );
  nand2_1 U29082 ( .ip1(\LUT[36][1] ), .ip2(n27477), .op(n25079) );
  nand2_1 U29083 ( .ip1(n27478), .ip2(\LUT[37][1] ), .op(n25078) );
  nand2_1 U29084 ( .ip1(n27479), .ip2(\LUT[32][1] ), .op(n25077) );
  nand3_1 U29085 ( .ip1(n25079), .ip2(n25078), .ip3(n25077), .op(n25080) );
  not_ab_or_c_or_d U29086 ( .ip1(n27485), .ip2(\LUT[40][1] ), .ip3(n25081), 
        .ip4(n25080), .op(n25085) );
  nand2_1 U29087 ( .ip1(n27487), .ip2(\LUT[35][1] ), .op(n25084) );
  nand2_1 U29088 ( .ip1(n27488), .ip2(\LUT[33][1] ), .op(n25083) );
  nand2_1 U29089 ( .ip1(n27486), .ip2(\LUT[34][1] ), .op(n25082) );
  nand4_1 U29090 ( .ip1(n25085), .ip2(n25084), .ip3(n25083), .ip4(n25082), 
        .op(n25086) );
  not_ab_or_c_or_d U29091 ( .ip1(n27495), .ip2(\LUT[29][1] ), .ip3(n25087), 
        .ip4(n25086), .op(n25088) );
  nor2_1 U29092 ( .ip1(n25088), .ip2(n27496), .op(n25107) );
  nand2_1 U29093 ( .ip1(n27498), .ip2(\LUT[48][1] ), .op(n25092) );
  nand2_1 U29094 ( .ip1(n27499), .ip2(\LUT[49][1] ), .op(n25091) );
  nand2_1 U29095 ( .ip1(n27500), .ip2(\LUT[53][1] ), .op(n25090) );
  nand2_1 U29096 ( .ip1(n27501), .ip2(\LUT[52][1] ), .op(n25089) );
  nand4_1 U29097 ( .ip1(n25092), .ip2(n25091), .ip3(n25090), .ip4(n25089), 
        .op(n25104) );
  and2_1 U29098 ( .ip1(n27520), .ip2(\LUT[47][1] ), .op(n25098) );
  nand2_1 U29099 ( .ip1(n27507), .ip2(\LUT[54][1] ), .op(n25096) );
  nand2_1 U29100 ( .ip1(n27508), .ip2(\LUT[55][1] ), .op(n25095) );
  nand2_1 U29101 ( .ip1(n27509), .ip2(\LUT[56][1] ), .op(n25094) );
  nand2_1 U29102 ( .ip1(n27510), .ip2(\LUT[51][1] ), .op(n25093) );
  nand4_1 U29103 ( .ip1(n25096), .ip2(n25095), .ip3(n25094), .ip4(n25093), 
        .op(n25097) );
  not_ab_or_c_or_d U29104 ( .ip1(n27517), .ip2(\LUT[50][1] ), .ip3(n25098), 
        .ip4(n25097), .op(n25102) );
  nand2_1 U29105 ( .ip1(n27518), .ip2(\LUT[44][1] ), .op(n25101) );
  nand2_1 U29106 ( .ip1(n27519), .ip2(\LUT[43][1] ), .op(n25100) );
  nand2_1 U29107 ( .ip1(n27506), .ip2(\LUT[45][1] ), .op(n25099) );
  nand4_1 U29108 ( .ip1(n25102), .ip2(n25101), .ip3(n25100), .ip4(n25099), 
        .op(n25103) );
  not_ab_or_c_or_d U29109 ( .ip1(n27527), .ip2(\LUT[46][1] ), .ip3(n25104), 
        .ip4(n25103), .op(n25105) );
  nor2_1 U29110 ( .ip1(n25105), .ip2(n27528), .op(n25106) );
  not_ab_or_c_or_d U29111 ( .ip1(n27533), .ip2(n25108), .ip3(n25107), .ip4(
        n25106), .op(n25109) );
  or2_1 U29112 ( .ip1(n25109), .ip2(n27265), .op(n25110) );
  nand2_1 U29113 ( .ip1(n25111), .ip2(n25110), .op(n25125) );
  nand2_1 U29114 ( .ip1(n27391), .ip2(\LUT[75][1] ), .op(n25123) );
  nand2_1 U29115 ( .ip1(n27373), .ip2(\LUT[82][1] ), .op(n25115) );
  nand2_1 U29116 ( .ip1(n27374), .ip2(\LUT[81][1] ), .op(n25114) );
  nand2_1 U29117 ( .ip1(n27375), .ip2(\LUT[84][1] ), .op(n25113) );
  nand2_1 U29118 ( .ip1(n27376), .ip2(\LUT[83][1] ), .op(n25112) );
  nand4_1 U29119 ( .ip1(n25115), .ip2(n25114), .ip3(n25113), .ip4(n25112), 
        .op(n25120) );
  nand2_1 U29120 ( .ip1(n27381), .ip2(\LUT[78][1] ), .op(n25118) );
  nand2_1 U29121 ( .ip1(n27382), .ip2(\LUT[79][1] ), .op(n25117) );
  nand2_1 U29122 ( .ip1(n27383), .ip2(\LUT[77][1] ), .op(n25116) );
  nand3_1 U29123 ( .ip1(n25118), .ip2(n25117), .ip3(n25116), .op(n25119) );
  not_ab_or_c_or_d U29124 ( .ip1(n27389), .ip2(\LUT[80][1] ), .ip3(n25120), 
        .ip4(n25119), .op(n25122) );
  nand2_1 U29125 ( .ip1(n27392), .ip2(\LUT[74][1] ), .op(n25121) );
  nand3_1 U29126 ( .ip1(n25123), .ip2(n25122), .ip3(n25121), .op(n25124) );
  not_ab_or_c_or_d U29127 ( .ip1(n27390), .ip2(\LUT[76][1] ), .ip3(n25125), 
        .ip4(n25124), .op(n25129) );
  nand2_1 U29128 ( .ip1(n27576), .ip2(\LUT[71][1] ), .op(n25128) );
  nand2_1 U29129 ( .ip1(n27569), .ip2(\LUT[73][1] ), .op(n25127) );
  nand2_1 U29130 ( .ip1(n27570), .ip2(\LUT[72][1] ), .op(n25126) );
  nand4_1 U29131 ( .ip1(n25129), .ip2(n25128), .ip3(n25127), .ip4(n25126), 
        .op(n25130) );
  nand2_1 U29132 ( .ip1(n27288), .ip2(n25130), .op(n25133) );
  nand2_1 U29133 ( .ip1(n27172), .ip2(\LUT[111][1] ), .op(n25132) );
  nand2_1 U29134 ( .ip1(n27165), .ip2(\LUT[108][1] ), .op(n25131) );
  nand4_1 U29135 ( .ip1(n25134), .ip2(n25133), .ip3(n25132), .ip4(n25131), 
        .op(n25135) );
  nand2_1 U29136 ( .ip1(n27589), .ip2(n25135), .op(n25137) );
  nand2_1 U29137 ( .ip1(sig_out[1]), .ip2(n27590), .op(n25136) );
  nand2_1 U29138 ( .ip1(n25137), .ip2(n25136), .op(n13464) );
  nand2_1 U29139 ( .ip1(n27333), .ip2(\LUT[95][2] ), .op(n25141) );
  nand2_1 U29140 ( .ip1(n27334), .ip2(\LUT[94][2] ), .op(n25140) );
  nand2_1 U29141 ( .ip1(n27335), .ip2(\LUT[98][2] ), .op(n25139) );
  nand2_1 U29142 ( .ip1(n27336), .ip2(\LUT[97][2] ), .op(n25138) );
  nand4_1 U29143 ( .ip1(n25141), .ip2(n25140), .ip3(n25139), .ip4(n25138), 
        .op(n25146) );
  nand2_1 U29144 ( .ip1(n27341), .ip2(\LUT[93][2] ), .op(n25144) );
  nand2_1 U29145 ( .ip1(n27342), .ip2(\LUT[92][2] ), .op(n25143) );
  nand2_1 U29146 ( .ip1(n27343), .ip2(\LUT[91][2] ), .op(n25142) );
  nand3_1 U29147 ( .ip1(n25144), .ip2(n25143), .ip3(n25142), .op(n25145) );
  not_ab_or_c_or_d U29148 ( .ip1(n27349), .ip2(\LUT[96][2] ), .ip3(n25146), 
        .ip4(n25145), .op(n25150) );
  nand2_1 U29149 ( .ip1(n27350), .ip2(\LUT[89][2] ), .op(n25149) );
  nand2_1 U29150 ( .ip1(n27351), .ip2(\LUT[90][2] ), .op(n25148) );
  nand2_1 U29151 ( .ip1(n27352), .ip2(\LUT[88][2] ), .op(n25147) );
  nand4_1 U29152 ( .ip1(n25150), .ip2(n25149), .ip3(n25148), .ip4(n25147), 
        .op(n25154) );
  nand2_1 U29153 ( .ip1(\LUT[85][2] ), .ip2(n27357), .op(n25152) );
  nand2_1 U29154 ( .ip1(\LUT[86][2] ), .ip2(n27358), .op(n25151) );
  nand2_1 U29155 ( .ip1(n25152), .ip2(n25151), .op(n25153) );
  not_ab_or_c_or_d U29156 ( .ip1(n27363), .ip2(\LUT[87][2] ), .ip3(n25154), 
        .ip4(n25153), .op(n25155) );
  nor2_1 U29157 ( .ip1(n25155), .ip2(n27142), .op(n25167) );
  and2_1 U29158 ( .ip1(n27317), .ip2(\LUT[105][2] ), .op(n25161) );
  nand2_1 U29159 ( .ip1(n27318), .ip2(\LUT[107][2] ), .op(n25159) );
  nand2_1 U29160 ( .ip1(n27319), .ip2(\LUT[104][2] ), .op(n25158) );
  nand2_1 U29161 ( .ip1(n27325), .ip2(\LUT[110][2] ), .op(n25157) );
  nand2_1 U29162 ( .ip1(n27309), .ip2(\LUT[109][2] ), .op(n25156) );
  nand4_1 U29163 ( .ip1(n25159), .ip2(n25158), .ip3(n25157), .ip4(n25156), 
        .op(n25160) );
  not_ab_or_c_or_d U29164 ( .ip1(\LUT[102][2] ), .ip2(n27326), .ip3(n25161), 
        .ip4(n25160), .op(n25165) );
  nand2_1 U29165 ( .ip1(n27370), .ip2(\LUT[100][2] ), .op(n25164) );
  nand2_1 U29166 ( .ip1(n27328), .ip2(\LUT[101][2] ), .op(n25163) );
  nand2_1 U29167 ( .ip1(n27327), .ip2(\LUT[103][2] ), .op(n25162) );
  nand4_1 U29168 ( .ip1(n25165), .ip2(n25164), .ip3(n25163), .ip4(n25162), 
        .op(n25166) );
  not_ab_or_c_or_d U29169 ( .ip1(\LUT[99][2] ), .ip2(n27156), .ip3(n25167), 
        .ip4(n25166), .op(n25168) );
  nor2_1 U29170 ( .ip1(n25168), .ip2(n27371), .op(n25181) );
  nand2_1 U29171 ( .ip1(n27582), .ip2(\LUT[115][2] ), .op(n25172) );
  nand2_1 U29172 ( .ip1(n27298), .ip2(\LUT[117][2] ), .op(n25171) );
  nand2_1 U29173 ( .ip1(n27299), .ip2(\LUT[118][2] ), .op(n25170) );
  nand2_1 U29174 ( .ip1(n27300), .ip2(\LUT[119][2] ), .op(n25169) );
  nand4_1 U29175 ( .ip1(n25172), .ip2(n25171), .ip3(n25170), .ip4(n25169), 
        .op(n25173) );
  or2_1 U29176 ( .ip1(n27297), .ip2(n25173), .op(n25175) );
  or2_1 U29177 ( .ip1(\LUT[116][2] ), .ip2(n25173), .op(n25174) );
  nand2_1 U29178 ( .ip1(n25175), .ip2(n25174), .op(n25179) );
  nand2_1 U29179 ( .ip1(n27583), .ip2(\LUT[113][2] ), .op(n25178) );
  nand2_1 U29180 ( .ip1(n27172), .ip2(\LUT[111][2] ), .op(n25177) );
  nand2_1 U29181 ( .ip1(n27305), .ip2(\LUT[114][2] ), .op(n25176) );
  nand4_1 U29182 ( .ip1(n25179), .ip2(n25178), .ip3(n25177), .ip4(n25176), 
        .op(n25180) );
  not_ab_or_c_or_d U29183 ( .ip1(n27581), .ip2(\LUT[106][2] ), .ip3(n25181), 
        .ip4(n25180), .op(n25299) );
  and2_1 U29184 ( .ip1(n27534), .ip2(\LUT[65][2] ), .op(n25187) );
  nand2_1 U29185 ( .ip1(n27548), .ip2(\LUT[67][2] ), .op(n25185) );
  nand2_1 U29186 ( .ip1(n27535), .ip2(\LUT[69][2] ), .op(n25184) );
  nand2_1 U29187 ( .ip1(n27536), .ip2(\LUT[70][2] ), .op(n25183) );
  nand2_1 U29188 ( .ip1(n27537), .ip2(\LUT[68][2] ), .op(n25182) );
  nand4_1 U29189 ( .ip1(n25185), .ip2(n25184), .ip3(n25183), .ip4(n25182), 
        .op(n25186) );
  not_ab_or_c_or_d U29190 ( .ip1(n27542), .ip2(\LUT[66][2] ), .ip3(n25187), 
        .ip4(n25186), .op(n25191) );
  nand2_1 U29191 ( .ip1(n27547), .ip2(\LUT[64][2] ), .op(n25190) );
  nand2_1 U29192 ( .ip1(n27556), .ip2(\LUT[63][2] ), .op(n25189) );
  nand2_1 U29193 ( .ip1(n27546), .ip2(\LUT[59][2] ), .op(n25188) );
  nand4_1 U29194 ( .ip1(n25191), .ip2(n25190), .ip3(n25189), .ip4(n25188), 
        .op(n25197) );
  nand2_1 U29195 ( .ip1(n27397), .ip2(\LUT[58][2] ), .op(n25195) );
  nand2_1 U29196 ( .ip1(n27563), .ip2(\LUT[62][2] ), .op(n25194) );
  nand2_1 U29197 ( .ip1(n27555), .ip2(\LUT[61][2] ), .op(n25193) );
  nand2_1 U29198 ( .ip1(n27554), .ip2(\LUT[60][2] ), .op(n25192) );
  nand4_1 U29199 ( .ip1(n25195), .ip2(n25194), .ip3(n25193), .ip4(n25192), 
        .op(n25196) );
  not_ab_or_c_or_d U29200 ( .ip1(n27553), .ip2(\LUT[57][2] ), .ip3(n25197), 
        .ip4(n25196), .op(n25198) );
  or2_1 U29201 ( .ip1(n25198), .ip2(n27265), .op(n25276) );
  nand2_1 U29202 ( .ip1(\LUT[27][2] ), .ip2(n27398), .op(n25201) );
  nand2_1 U29203 ( .ip1(n27405), .ip2(\LUT[25][2] ), .op(n25200) );
  nand2_1 U29204 ( .ip1(n27400), .ip2(\LUT[28][2] ), .op(n25199) );
  nand3_1 U29205 ( .ip1(n25201), .ip2(n25200), .ip3(n25199), .op(n25206) );
  nand2_1 U29206 ( .ip1(\LUT[24][2] ), .ip2(n27404), .op(n25204) );
  nand2_1 U29207 ( .ip1(n27406), .ip2(\LUT[23][2] ), .op(n25203) );
  nand2_1 U29208 ( .ip1(n27399), .ip2(\LUT[26][2] ), .op(n25202) );
  nand3_1 U29209 ( .ip1(n25204), .ip2(n25203), .ip3(n25202), .op(n25205) );
  not_ab_or_c_or_d U29210 ( .ip1(n27460), .ip2(\LUT[19][2] ), .ip3(n25206), 
        .ip4(n25205), .op(n25235) );
  nand2_1 U29211 ( .ip1(\LUT[2][2] ), .ip2(n27413), .op(n25208) );
  nand2_1 U29212 ( .ip1(\LUT[3][2] ), .ip2(n27414), .op(n25207) );
  nand2_1 U29213 ( .ip1(n25208), .ip2(n25207), .op(n25224) );
  nand2_1 U29214 ( .ip1(n27427), .ip2(\LUT[12][2] ), .op(n25212) );
  nand2_1 U29215 ( .ip1(n27417), .ip2(\LUT[7][2] ), .op(n25211) );
  nand2_1 U29216 ( .ip1(n27420), .ip2(\LUT[13][2] ), .op(n25210) );
  nand2_1 U29217 ( .ip1(n27419), .ip2(\LUT[14][2] ), .op(n25209) );
  nand4_1 U29218 ( .ip1(n25212), .ip2(n25211), .ip3(n25210), .ip4(n25209), 
        .op(n25218) );
  nand2_1 U29219 ( .ip1(n27425), .ip2(\LUT[10][2] ), .op(n25216) );
  nand2_1 U29220 ( .ip1(n27428), .ip2(\LUT[6][2] ), .op(n25215) );
  nand2_1 U29221 ( .ip1(n27426), .ip2(\LUT[8][2] ), .op(n25214) );
  nand2_1 U29222 ( .ip1(n27435), .ip2(\LUT[11][2] ), .op(n25213) );
  nand4_1 U29223 ( .ip1(n25216), .ip2(n25215), .ip3(n25214), .ip4(n25213), 
        .op(n25217) );
  not_ab_or_c_or_d U29224 ( .ip1(n27418), .ip2(\LUT[9][2] ), .ip3(n25218), 
        .ip4(n25217), .op(n25222) );
  nand2_1 U29225 ( .ip1(n27445), .ip2(\LUT[1][2] ), .op(n25221) );
  nand2_1 U29226 ( .ip1(n27437), .ip2(\LUT[4][2] ), .op(n25220) );
  nand2_1 U29227 ( .ip1(n27438), .ip2(\LUT[5][2] ), .op(n25219) );
  nand4_1 U29228 ( .ip1(n25222), .ip2(n25221), .ip3(n25220), .ip4(n25219), 
        .op(n25223) );
  not_ab_or_c_or_d U29229 ( .ip1(n27436), .ip2(\LUT[0][2] ), .ip3(n25224), 
        .ip4(n25223), .op(n25225) );
  nor2_1 U29230 ( .ip1(n25225), .ip2(n27446), .op(n25231) );
  nand2_1 U29231 ( .ip1(n27450), .ip2(\LUT[21][2] ), .op(n25229) );
  nand2_1 U29232 ( .ip1(n27451), .ip2(\LUT[16][2] ), .op(n25228) );
  nand2_1 U29233 ( .ip1(n27448), .ip2(\LUT[18][2] ), .op(n25227) );
  nand2_1 U29234 ( .ip1(n27449), .ip2(\LUT[20][2] ), .op(n25226) );
  nand4_1 U29235 ( .ip1(n25229), .ip2(n25228), .ip3(n25227), .ip4(n25226), 
        .op(n25230) );
  not_ab_or_c_or_d U29236 ( .ip1(\LUT[15][2] ), .ip2(n27458), .ip3(n25231), 
        .ip4(n25230), .op(n25234) );
  nand2_1 U29237 ( .ip1(n27459), .ip2(\LUT[17][2] ), .op(n25233) );
  nand2_1 U29238 ( .ip1(n27412), .ip2(\LUT[22][2] ), .op(n25232) );
  nand4_1 U29239 ( .ip1(n25235), .ip2(n25234), .ip3(n25233), .ip4(n25232), 
        .op(n25273) );
  nand2_1 U29240 ( .ip1(n27498), .ip2(\LUT[48][2] ), .op(n25239) );
  nand2_1 U29241 ( .ip1(n27499), .ip2(\LUT[49][2] ), .op(n25238) );
  nand2_1 U29242 ( .ip1(n27500), .ip2(\LUT[53][2] ), .op(n25237) );
  nand2_1 U29243 ( .ip1(n27501), .ip2(\LUT[52][2] ), .op(n25236) );
  nand4_1 U29244 ( .ip1(n25239), .ip2(n25238), .ip3(n25237), .ip4(n25236), 
        .op(n25251) );
  and2_1 U29245 ( .ip1(n27518), .ip2(\LUT[44][2] ), .op(n25245) );
  nand2_1 U29246 ( .ip1(n27507), .ip2(\LUT[54][2] ), .op(n25243) );
  nand2_1 U29247 ( .ip1(n27509), .ip2(\LUT[56][2] ), .op(n25242) );
  nand2_1 U29248 ( .ip1(n27508), .ip2(\LUT[55][2] ), .op(n25241) );
  nand2_1 U29249 ( .ip1(n27510), .ip2(\LUT[51][2] ), .op(n25240) );
  nand4_1 U29250 ( .ip1(n25243), .ip2(n25242), .ip3(n25241), .ip4(n25240), 
        .op(n25244) );
  not_ab_or_c_or_d U29251 ( .ip1(n27517), .ip2(\LUT[50][2] ), .ip3(n25245), 
        .ip4(n25244), .op(n25249) );
  nand2_1 U29252 ( .ip1(n27506), .ip2(\LUT[45][2] ), .op(n25248) );
  nand2_1 U29253 ( .ip1(n27519), .ip2(\LUT[43][2] ), .op(n25247) );
  nand2_1 U29254 ( .ip1(n27520), .ip2(\LUT[47][2] ), .op(n25246) );
  nand4_1 U29255 ( .ip1(n25249), .ip2(n25248), .ip3(n25247), .ip4(n25246), 
        .op(n25250) );
  not_ab_or_c_or_d U29256 ( .ip1(n27527), .ip2(\LUT[46][2] ), .ip3(n25251), 
        .ip4(n25250), .op(n25252) );
  nor2_1 U29257 ( .ip1(n25252), .ip2(n27528), .op(n25272) );
  nand2_1 U29258 ( .ip1(\LUT[31][2] ), .ip2(n27465), .op(n25254) );
  nand2_1 U29259 ( .ip1(\LUT[30][2] ), .ip2(n27466), .op(n25253) );
  nand2_1 U29260 ( .ip1(n25254), .ip2(n25253), .op(n25269) );
  nand2_1 U29261 ( .ip1(n27470), .ip2(\LUT[38][2] ), .op(n25258) );
  nand2_1 U29262 ( .ip1(n27469), .ip2(\LUT[39][2] ), .op(n25257) );
  nand2_1 U29263 ( .ip1(n27471), .ip2(\LUT[41][2] ), .op(n25256) );
  nand2_1 U29264 ( .ip1(n27472), .ip2(\LUT[42][2] ), .op(n25255) );
  nand4_1 U29265 ( .ip1(n25258), .ip2(n25257), .ip3(n25256), .ip4(n25255), 
        .op(n25263) );
  nand2_1 U29266 ( .ip1(\LUT[36][2] ), .ip2(n27477), .op(n25261) );
  nand2_1 U29267 ( .ip1(n27479), .ip2(\LUT[32][2] ), .op(n25260) );
  nand2_1 U29268 ( .ip1(n27478), .ip2(\LUT[37][2] ), .op(n25259) );
  nand3_1 U29269 ( .ip1(n25261), .ip2(n25260), .ip3(n25259), .op(n25262) );
  not_ab_or_c_or_d U29270 ( .ip1(n27485), .ip2(\LUT[40][2] ), .ip3(n25263), 
        .ip4(n25262), .op(n25267) );
  nand2_1 U29271 ( .ip1(n27486), .ip2(\LUT[34][2] ), .op(n25266) );
  nand2_1 U29272 ( .ip1(n27488), .ip2(\LUT[33][2] ), .op(n25265) );
  nand2_1 U29273 ( .ip1(n27487), .ip2(\LUT[35][2] ), .op(n25264) );
  nand4_1 U29274 ( .ip1(n25267), .ip2(n25266), .ip3(n25265), .ip4(n25264), 
        .op(n25268) );
  not_ab_or_c_or_d U29275 ( .ip1(n27495), .ip2(\LUT[29][2] ), .ip3(n25269), 
        .ip4(n25268), .op(n25270) );
  nor2_1 U29276 ( .ip1(n25270), .ip2(n27496), .op(n25271) );
  not_ab_or_c_or_d U29277 ( .ip1(n27533), .ip2(n25273), .ip3(n25272), .ip4(
        n25271), .op(n25274) );
  or2_1 U29278 ( .ip1(n25274), .ip2(n27265), .op(n25275) );
  nand2_1 U29279 ( .ip1(n25276), .ip2(n25275), .op(n25290) );
  nand2_1 U29280 ( .ip1(n27391), .ip2(\LUT[75][2] ), .op(n25288) );
  nand2_1 U29281 ( .ip1(n27373), .ip2(\LUT[82][2] ), .op(n25280) );
  nand2_1 U29282 ( .ip1(n27374), .ip2(\LUT[81][2] ), .op(n25279) );
  nand2_1 U29283 ( .ip1(n27375), .ip2(\LUT[84][2] ), .op(n25278) );
  nand2_1 U29284 ( .ip1(n27376), .ip2(\LUT[83][2] ), .op(n25277) );
  nand4_1 U29285 ( .ip1(n25280), .ip2(n25279), .ip3(n25278), .ip4(n25277), 
        .op(n25285) );
  nand2_1 U29286 ( .ip1(\LUT[78][2] ), .ip2(n27381), .op(n25283) );
  nand2_1 U29287 ( .ip1(n27382), .ip2(\LUT[79][2] ), .op(n25282) );
  nand2_1 U29288 ( .ip1(n27383), .ip2(\LUT[77][2] ), .op(n25281) );
  nand3_1 U29289 ( .ip1(n25283), .ip2(n25282), .ip3(n25281), .op(n25284) );
  not_ab_or_c_or_d U29290 ( .ip1(n27389), .ip2(\LUT[80][2] ), .ip3(n25285), 
        .ip4(n25284), .op(n25287) );
  nand2_1 U29291 ( .ip1(n27392), .ip2(\LUT[74][2] ), .op(n25286) );
  nand3_1 U29292 ( .ip1(n25288), .ip2(n25287), .ip3(n25286), .op(n25289) );
  not_ab_or_c_or_d U29293 ( .ip1(n27390), .ip2(\LUT[76][2] ), .ip3(n25290), 
        .ip4(n25289), .op(n25294) );
  nand2_1 U29294 ( .ip1(n27576), .ip2(\LUT[71][2] ), .op(n25293) );
  nand2_1 U29295 ( .ip1(n27569), .ip2(\LUT[73][2] ), .op(n25292) );
  nand2_1 U29296 ( .ip1(n27570), .ip2(\LUT[72][2] ), .op(n25291) );
  nand4_1 U29297 ( .ip1(n25294), .ip2(n25293), .ip3(n25292), .ip4(n25291), 
        .op(n25295) );
  nand2_1 U29298 ( .ip1(n27288), .ip2(n25295), .op(n25298) );
  nand2_1 U29299 ( .ip1(n27289), .ip2(\LUT[112][2] ), .op(n25297) );
  nand2_1 U29300 ( .ip1(n27165), .ip2(\LUT[108][2] ), .op(n25296) );
  nand4_1 U29301 ( .ip1(n25299), .ip2(n25298), .ip3(n25297), .ip4(n25296), 
        .op(n25300) );
  nand2_1 U29302 ( .ip1(n27589), .ip2(n25300), .op(n25302) );
  nand2_1 U29303 ( .ip1(sig_out[2]), .ip2(n27590), .op(n25301) );
  nand2_1 U29304 ( .ip1(n25302), .ip2(n25301), .op(n13463) );
  nand2_1 U29305 ( .ip1(n27333), .ip2(\LUT[95][3] ), .op(n25306) );
  nand2_1 U29306 ( .ip1(n27334), .ip2(\LUT[94][3] ), .op(n25305) );
  nand2_1 U29307 ( .ip1(n27336), .ip2(\LUT[97][3] ), .op(n25304) );
  nand2_1 U29308 ( .ip1(n27335), .ip2(\LUT[98][3] ), .op(n25303) );
  nand4_1 U29309 ( .ip1(n25306), .ip2(n25305), .ip3(n25304), .ip4(n25303), 
        .op(n25311) );
  nand2_1 U29310 ( .ip1(n27341), .ip2(\LUT[93][3] ), .op(n25309) );
  nand2_1 U29311 ( .ip1(n27342), .ip2(\LUT[92][3] ), .op(n25308) );
  nand2_1 U29312 ( .ip1(n27343), .ip2(\LUT[91][3] ), .op(n25307) );
  nand3_1 U29313 ( .ip1(n25309), .ip2(n25308), .ip3(n25307), .op(n25310) );
  not_ab_or_c_or_d U29314 ( .ip1(n27349), .ip2(\LUT[96][3] ), .ip3(n25311), 
        .ip4(n25310), .op(n25315) );
  nand2_1 U29315 ( .ip1(n27350), .ip2(\LUT[89][3] ), .op(n25314) );
  nand2_1 U29316 ( .ip1(n27351), .ip2(\LUT[90][3] ), .op(n25313) );
  nand2_1 U29317 ( .ip1(n27352), .ip2(\LUT[88][3] ), .op(n25312) );
  nand4_1 U29318 ( .ip1(n25315), .ip2(n25314), .ip3(n25313), .ip4(n25312), 
        .op(n25319) );
  nand2_1 U29319 ( .ip1(\LUT[85][3] ), .ip2(n27357), .op(n25317) );
  nand2_1 U29320 ( .ip1(\LUT[86][3] ), .ip2(n27358), .op(n25316) );
  nand2_1 U29321 ( .ip1(n25317), .ip2(n25316), .op(n25318) );
  not_ab_or_c_or_d U29322 ( .ip1(n27363), .ip2(\LUT[87][3] ), .ip3(n25319), 
        .ip4(n25318), .op(n25320) );
  nor2_1 U29323 ( .ip1(n25320), .ip2(n27142), .op(n25332) );
  and2_1 U29324 ( .ip1(n27317), .ip2(\LUT[105][3] ), .op(n25326) );
  nand2_1 U29325 ( .ip1(n27318), .ip2(\LUT[107][3] ), .op(n25324) );
  nand2_1 U29326 ( .ip1(n27319), .ip2(\LUT[104][3] ), .op(n25323) );
  nand2_1 U29327 ( .ip1(n27325), .ip2(\LUT[110][3] ), .op(n25322) );
  nand2_1 U29328 ( .ip1(n27309), .ip2(\LUT[109][3] ), .op(n25321) );
  nand4_1 U29329 ( .ip1(n25324), .ip2(n25323), .ip3(n25322), .ip4(n25321), 
        .op(n25325) );
  not_ab_or_c_or_d U29330 ( .ip1(\LUT[102][3] ), .ip2(n27326), .ip3(n25326), 
        .ip4(n25325), .op(n25330) );
  nand2_1 U29331 ( .ip1(n27370), .ip2(\LUT[100][3] ), .op(n25329) );
  nand2_1 U29332 ( .ip1(n27328), .ip2(\LUT[101][3] ), .op(n25328) );
  nand2_1 U29333 ( .ip1(n27327), .ip2(\LUT[103][3] ), .op(n25327) );
  nand4_1 U29334 ( .ip1(n25330), .ip2(n25329), .ip3(n25328), .ip4(n25327), 
        .op(n25331) );
  not_ab_or_c_or_d U29335 ( .ip1(\LUT[99][3] ), .ip2(n27156), .ip3(n25332), 
        .ip4(n25331), .op(n25333) );
  nor2_1 U29336 ( .ip1(n25333), .ip2(n27371), .op(n25346) );
  nand2_1 U29337 ( .ip1(n27582), .ip2(\LUT[115][3] ), .op(n25337) );
  nand2_1 U29338 ( .ip1(n27298), .ip2(\LUT[117][3] ), .op(n25336) );
  nand2_1 U29339 ( .ip1(n27299), .ip2(\LUT[118][3] ), .op(n25335) );
  nand2_1 U29340 ( .ip1(n27300), .ip2(\LUT[119][3] ), .op(n25334) );
  nand4_1 U29341 ( .ip1(n25337), .ip2(n25336), .ip3(n25335), .ip4(n25334), 
        .op(n25338) );
  or2_1 U29342 ( .ip1(n27297), .ip2(n25338), .op(n25340) );
  or2_1 U29343 ( .ip1(\LUT[116][3] ), .ip2(n25338), .op(n25339) );
  nand2_1 U29344 ( .ip1(n25340), .ip2(n25339), .op(n25344) );
  nand2_1 U29345 ( .ip1(n27583), .ip2(\LUT[113][3] ), .op(n25343) );
  nand2_1 U29346 ( .ip1(n27172), .ip2(\LUT[111][3] ), .op(n25342) );
  nand2_1 U29347 ( .ip1(n27305), .ip2(\LUT[114][3] ), .op(n25341) );
  nand4_1 U29348 ( .ip1(n25344), .ip2(n25343), .ip3(n25342), .ip4(n25341), 
        .op(n25345) );
  not_ab_or_c_or_d U29349 ( .ip1(n27581), .ip2(\LUT[106][3] ), .ip3(n25346), 
        .ip4(n25345), .op(n25464) );
  and2_1 U29350 ( .ip1(n27534), .ip2(\LUT[65][3] ), .op(n25352) );
  nand2_1 U29351 ( .ip1(n27548), .ip2(\LUT[67][3] ), .op(n25350) );
  nand2_1 U29352 ( .ip1(n27536), .ip2(\LUT[70][3] ), .op(n25349) );
  nand2_1 U29353 ( .ip1(n27535), .ip2(\LUT[69][3] ), .op(n25348) );
  nand2_1 U29354 ( .ip1(n27537), .ip2(\LUT[68][3] ), .op(n25347) );
  nand4_1 U29355 ( .ip1(n25350), .ip2(n25349), .ip3(n25348), .ip4(n25347), 
        .op(n25351) );
  not_ab_or_c_or_d U29356 ( .ip1(n27542), .ip2(\LUT[66][3] ), .ip3(n25352), 
        .ip4(n25351), .op(n25356) );
  nand2_1 U29357 ( .ip1(n27547), .ip2(\LUT[64][3] ), .op(n25355) );
  nand2_1 U29358 ( .ip1(n27563), .ip2(\LUT[62][3] ), .op(n25354) );
  nand2_1 U29359 ( .ip1(n27546), .ip2(\LUT[59][3] ), .op(n25353) );
  nand4_1 U29360 ( .ip1(n25356), .ip2(n25355), .ip3(n25354), .ip4(n25353), 
        .op(n25362) );
  nand2_1 U29361 ( .ip1(n27397), .ip2(\LUT[58][3] ), .op(n25360) );
  nand2_1 U29362 ( .ip1(n27554), .ip2(\LUT[60][3] ), .op(n25359) );
  nand2_1 U29363 ( .ip1(n27556), .ip2(\LUT[63][3] ), .op(n25358) );
  nand2_1 U29364 ( .ip1(n27555), .ip2(\LUT[61][3] ), .op(n25357) );
  nand4_1 U29365 ( .ip1(n25360), .ip2(n25359), .ip3(n25358), .ip4(n25357), 
        .op(n25361) );
  not_ab_or_c_or_d U29366 ( .ip1(n27553), .ip2(\LUT[57][3] ), .ip3(n25362), 
        .ip4(n25361), .op(n25363) );
  or2_1 U29367 ( .ip1(n25363), .ip2(n27265), .op(n25441) );
  nand2_1 U29368 ( .ip1(\LUT[27][3] ), .ip2(n27398), .op(n25366) );
  nand2_1 U29369 ( .ip1(n27405), .ip2(\LUT[25][3] ), .op(n25365) );
  nand2_1 U29370 ( .ip1(n27400), .ip2(\LUT[28][3] ), .op(n25364) );
  nand3_1 U29371 ( .ip1(n25366), .ip2(n25365), .ip3(n25364), .op(n25371) );
  nand2_1 U29372 ( .ip1(\LUT[24][3] ), .ip2(n27404), .op(n25369) );
  nand2_1 U29373 ( .ip1(n27399), .ip2(\LUT[26][3] ), .op(n25368) );
  nand2_1 U29374 ( .ip1(n27406), .ip2(\LUT[23][3] ), .op(n25367) );
  nand3_1 U29375 ( .ip1(n25369), .ip2(n25368), .ip3(n25367), .op(n25370) );
  not_ab_or_c_or_d U29376 ( .ip1(n27460), .ip2(\LUT[19][3] ), .ip3(n25371), 
        .ip4(n25370), .op(n25400) );
  nand2_1 U29377 ( .ip1(\LUT[2][3] ), .ip2(n27413), .op(n25373) );
  nand2_1 U29378 ( .ip1(\LUT[3][3] ), .ip2(n27414), .op(n25372) );
  nand2_1 U29379 ( .ip1(n25373), .ip2(n25372), .op(n25389) );
  nand2_1 U29380 ( .ip1(n27418), .ip2(\LUT[9][3] ), .op(n25377) );
  nand2_1 U29381 ( .ip1(n27428), .ip2(\LUT[6][3] ), .op(n25376) );
  nand2_1 U29382 ( .ip1(n27420), .ip2(\LUT[13][3] ), .op(n25375) );
  nand2_1 U29383 ( .ip1(n27419), .ip2(\LUT[14][3] ), .op(n25374) );
  nand4_1 U29384 ( .ip1(n25377), .ip2(n25376), .ip3(n25375), .ip4(n25374), 
        .op(n25383) );
  nand2_1 U29385 ( .ip1(n27427), .ip2(\LUT[12][3] ), .op(n25381) );
  nand2_1 U29386 ( .ip1(n27425), .ip2(\LUT[10][3] ), .op(n25380) );
  nand2_1 U29387 ( .ip1(n27426), .ip2(\LUT[8][3] ), .op(n25379) );
  nand2_1 U29388 ( .ip1(n27417), .ip2(\LUT[7][3] ), .op(n25378) );
  nand4_1 U29389 ( .ip1(n25381), .ip2(n25380), .ip3(n25379), .ip4(n25378), 
        .op(n25382) );
  not_ab_or_c_or_d U29390 ( .ip1(n27435), .ip2(\LUT[11][3] ), .ip3(n25383), 
        .ip4(n25382), .op(n25387) );
  nand2_1 U29391 ( .ip1(n27436), .ip2(\LUT[0][3] ), .op(n25386) );
  nand2_1 U29392 ( .ip1(n27437), .ip2(\LUT[4][3] ), .op(n25385) );
  nand2_1 U29393 ( .ip1(n27438), .ip2(\LUT[5][3] ), .op(n25384) );
  nand4_1 U29394 ( .ip1(n25387), .ip2(n25386), .ip3(n25385), .ip4(n25384), 
        .op(n25388) );
  not_ab_or_c_or_d U29395 ( .ip1(n27445), .ip2(\LUT[1][3] ), .ip3(n25389), 
        .ip4(n25388), .op(n25390) );
  nor2_1 U29396 ( .ip1(n25390), .ip2(n27446), .op(n25396) );
  nand2_1 U29397 ( .ip1(n27451), .ip2(\LUT[16][3] ), .op(n25394) );
  nand2_1 U29398 ( .ip1(n27450), .ip2(\LUT[21][3] ), .op(n25393) );
  nand2_1 U29399 ( .ip1(n27448), .ip2(\LUT[18][3] ), .op(n25392) );
  nand2_1 U29400 ( .ip1(n27449), .ip2(\LUT[20][3] ), .op(n25391) );
  nand4_1 U29401 ( .ip1(n25394), .ip2(n25393), .ip3(n25392), .ip4(n25391), 
        .op(n25395) );
  not_ab_or_c_or_d U29402 ( .ip1(\LUT[15][3] ), .ip2(n27458), .ip3(n25396), 
        .ip4(n25395), .op(n25399) );
  nand2_1 U29403 ( .ip1(n27412), .ip2(\LUT[22][3] ), .op(n25398) );
  nand2_1 U29404 ( .ip1(n27459), .ip2(\LUT[17][3] ), .op(n25397) );
  nand4_1 U29405 ( .ip1(n25400), .ip2(n25399), .ip3(n25398), .ip4(n25397), 
        .op(n25438) );
  nand2_1 U29406 ( .ip1(n27499), .ip2(\LUT[49][3] ), .op(n25404) );
  nand2_1 U29407 ( .ip1(n27498), .ip2(\LUT[48][3] ), .op(n25403) );
  nand2_1 U29408 ( .ip1(n27500), .ip2(\LUT[53][3] ), .op(n25402) );
  nand2_1 U29409 ( .ip1(n27501), .ip2(\LUT[52][3] ), .op(n25401) );
  nand4_1 U29410 ( .ip1(n25404), .ip2(n25403), .ip3(n25402), .ip4(n25401), 
        .op(n25416) );
  and2_1 U29411 ( .ip1(n27520), .ip2(\LUT[47][3] ), .op(n25410) );
  nand2_1 U29412 ( .ip1(n27507), .ip2(\LUT[54][3] ), .op(n25408) );
  nand2_1 U29413 ( .ip1(n27508), .ip2(\LUT[55][3] ), .op(n25407) );
  nand2_1 U29414 ( .ip1(n27509), .ip2(\LUT[56][3] ), .op(n25406) );
  nand2_1 U29415 ( .ip1(n27510), .ip2(\LUT[51][3] ), .op(n25405) );
  nand4_1 U29416 ( .ip1(n25408), .ip2(n25407), .ip3(n25406), .ip4(n25405), 
        .op(n25409) );
  not_ab_or_c_or_d U29417 ( .ip1(n27517), .ip2(\LUT[50][3] ), .ip3(n25410), 
        .ip4(n25409), .op(n25414) );
  nand2_1 U29418 ( .ip1(n27518), .ip2(\LUT[44][3] ), .op(n25413) );
  nand2_1 U29419 ( .ip1(n27519), .ip2(\LUT[43][3] ), .op(n25412) );
  nand2_1 U29420 ( .ip1(n27506), .ip2(\LUT[45][3] ), .op(n25411) );
  nand4_1 U29421 ( .ip1(n25414), .ip2(n25413), .ip3(n25412), .ip4(n25411), 
        .op(n25415) );
  not_ab_or_c_or_d U29422 ( .ip1(n27527), .ip2(\LUT[46][3] ), .ip3(n25416), 
        .ip4(n25415), .op(n25417) );
  nor2_1 U29423 ( .ip1(n25417), .ip2(n27528), .op(n25437) );
  nand2_1 U29424 ( .ip1(\LUT[31][3] ), .ip2(n27465), .op(n25419) );
  nand2_1 U29425 ( .ip1(\LUT[30][3] ), .ip2(n27466), .op(n25418) );
  nand2_1 U29426 ( .ip1(n25419), .ip2(n25418), .op(n25434) );
  nand2_1 U29427 ( .ip1(n27469), .ip2(\LUT[39][3] ), .op(n25423) );
  nand2_1 U29428 ( .ip1(n27470), .ip2(\LUT[38][3] ), .op(n25422) );
  nand2_1 U29429 ( .ip1(n27471), .ip2(\LUT[41][3] ), .op(n25421) );
  nand2_1 U29430 ( .ip1(n27472), .ip2(\LUT[42][3] ), .op(n25420) );
  nand4_1 U29431 ( .ip1(n25423), .ip2(n25422), .ip3(n25421), .ip4(n25420), 
        .op(n25428) );
  nand2_1 U29432 ( .ip1(\LUT[36][3] ), .ip2(n27477), .op(n25426) );
  nand2_1 U29433 ( .ip1(n27478), .ip2(\LUT[37][3] ), .op(n25425) );
  nand2_1 U29434 ( .ip1(n27479), .ip2(\LUT[32][3] ), .op(n25424) );
  nand3_1 U29435 ( .ip1(n25426), .ip2(n25425), .ip3(n25424), .op(n25427) );
  not_ab_or_c_or_d U29436 ( .ip1(n27485), .ip2(\LUT[40][3] ), .ip3(n25428), 
        .ip4(n25427), .op(n25432) );
  nand2_1 U29437 ( .ip1(n27488), .ip2(\LUT[33][3] ), .op(n25431) );
  nand2_1 U29438 ( .ip1(n27486), .ip2(\LUT[34][3] ), .op(n25430) );
  nand2_1 U29439 ( .ip1(n27487), .ip2(\LUT[35][3] ), .op(n25429) );
  nand4_1 U29440 ( .ip1(n25432), .ip2(n25431), .ip3(n25430), .ip4(n25429), 
        .op(n25433) );
  not_ab_or_c_or_d U29441 ( .ip1(n27495), .ip2(\LUT[29][3] ), .ip3(n25434), 
        .ip4(n25433), .op(n25435) );
  nor2_1 U29442 ( .ip1(n25435), .ip2(n27496), .op(n25436) );
  not_ab_or_c_or_d U29443 ( .ip1(n27533), .ip2(n25438), .ip3(n25437), .ip4(
        n25436), .op(n25439) );
  or2_1 U29444 ( .ip1(n25439), .ip2(n27265), .op(n25440) );
  nand2_1 U29445 ( .ip1(n25441), .ip2(n25440), .op(n25455) );
  nand2_1 U29446 ( .ip1(n27391), .ip2(\LUT[75][3] ), .op(n25453) );
  nand2_1 U29447 ( .ip1(n27373), .ip2(\LUT[82][3] ), .op(n25445) );
  nand2_1 U29448 ( .ip1(n27374), .ip2(\LUT[81][3] ), .op(n25444) );
  nand2_1 U29449 ( .ip1(n27375), .ip2(\LUT[84][3] ), .op(n25443) );
  nand2_1 U29450 ( .ip1(n27376), .ip2(\LUT[83][3] ), .op(n25442) );
  nand4_1 U29451 ( .ip1(n25445), .ip2(n25444), .ip3(n25443), .ip4(n25442), 
        .op(n25450) );
  nand2_1 U29452 ( .ip1(\LUT[78][3] ), .ip2(n27381), .op(n25448) );
  nand2_1 U29453 ( .ip1(n27382), .ip2(\LUT[79][3] ), .op(n25447) );
  nand2_1 U29454 ( .ip1(n27383), .ip2(\LUT[77][3] ), .op(n25446) );
  nand3_1 U29455 ( .ip1(n25448), .ip2(n25447), .ip3(n25446), .op(n25449) );
  not_ab_or_c_or_d U29456 ( .ip1(n27389), .ip2(\LUT[80][3] ), .ip3(n25450), 
        .ip4(n25449), .op(n25452) );
  nand2_1 U29457 ( .ip1(n27392), .ip2(\LUT[74][3] ), .op(n25451) );
  nand3_1 U29458 ( .ip1(n25453), .ip2(n25452), .ip3(n25451), .op(n25454) );
  not_ab_or_c_or_d U29459 ( .ip1(n27390), .ip2(\LUT[76][3] ), .ip3(n25455), 
        .ip4(n25454), .op(n25459) );
  nand2_1 U29460 ( .ip1(n27576), .ip2(\LUT[71][3] ), .op(n25458) );
  nand2_1 U29461 ( .ip1(n27570), .ip2(\LUT[72][3] ), .op(n25457) );
  nand2_1 U29462 ( .ip1(n27569), .ip2(\LUT[73][3] ), .op(n25456) );
  nand4_1 U29463 ( .ip1(n25459), .ip2(n25458), .ip3(n25457), .ip4(n25456), 
        .op(n25460) );
  nand2_1 U29464 ( .ip1(n27288), .ip2(n25460), .op(n25463) );
  nand2_1 U29465 ( .ip1(n27165), .ip2(\LUT[108][3] ), .op(n25462) );
  nand2_1 U29466 ( .ip1(n27289), .ip2(\LUT[112][3] ), .op(n25461) );
  nand4_1 U29467 ( .ip1(n25464), .ip2(n25463), .ip3(n25462), .ip4(n25461), 
        .op(n25465) );
  nand2_1 U29468 ( .ip1(n27589), .ip2(n25465), .op(n25467) );
  nand2_1 U29469 ( .ip1(sig_out[3]), .ip2(n27590), .op(n25466) );
  nand2_1 U29470 ( .ip1(n25467), .ip2(n25466), .op(n13462) );
  nand2_1 U29471 ( .ip1(n27333), .ip2(\LUT[95][4] ), .op(n25471) );
  nand2_1 U29472 ( .ip1(n27334), .ip2(\LUT[94][4] ), .op(n25470) );
  nand2_1 U29473 ( .ip1(n27336), .ip2(\LUT[97][4] ), .op(n25469) );
  nand2_1 U29474 ( .ip1(n27335), .ip2(\LUT[98][4] ), .op(n25468) );
  nand4_1 U29475 ( .ip1(n25471), .ip2(n25470), .ip3(n25469), .ip4(n25468), 
        .op(n25476) );
  nand2_1 U29476 ( .ip1(n27341), .ip2(\LUT[93][4] ), .op(n25474) );
  nand2_1 U29477 ( .ip1(n27342), .ip2(\LUT[92][4] ), .op(n25473) );
  nand2_1 U29478 ( .ip1(n27343), .ip2(\LUT[91][4] ), .op(n25472) );
  nand3_1 U29479 ( .ip1(n25474), .ip2(n25473), .ip3(n25472), .op(n25475) );
  not_ab_or_c_or_d U29480 ( .ip1(n27349), .ip2(\LUT[96][4] ), .ip3(n25476), 
        .ip4(n25475), .op(n25480) );
  nand2_1 U29481 ( .ip1(n27350), .ip2(\LUT[89][4] ), .op(n25479) );
  nand2_1 U29482 ( .ip1(n27351), .ip2(\LUT[90][4] ), .op(n25478) );
  nand2_1 U29483 ( .ip1(n27352), .ip2(\LUT[88][4] ), .op(n25477) );
  nand4_1 U29484 ( .ip1(n25480), .ip2(n25479), .ip3(n25478), .ip4(n25477), 
        .op(n25484) );
  nand2_1 U29485 ( .ip1(\LUT[85][4] ), .ip2(n27357), .op(n25482) );
  nand2_1 U29486 ( .ip1(\LUT[86][4] ), .ip2(n27358), .op(n25481) );
  nand2_1 U29487 ( .ip1(n25482), .ip2(n25481), .op(n25483) );
  not_ab_or_c_or_d U29488 ( .ip1(n27363), .ip2(\LUT[87][4] ), .ip3(n25484), 
        .ip4(n25483), .op(n25485) );
  nor2_1 U29489 ( .ip1(n25485), .ip2(n27142), .op(n25497) );
  and2_1 U29490 ( .ip1(n27317), .ip2(\LUT[105][4] ), .op(n25491) );
  nand2_1 U29491 ( .ip1(n27318), .ip2(\LUT[107][4] ), .op(n25489) );
  nand2_1 U29492 ( .ip1(n27319), .ip2(\LUT[104][4] ), .op(n25488) );
  nand2_1 U29493 ( .ip1(n27309), .ip2(\LUT[109][4] ), .op(n25487) );
  nand2_1 U29494 ( .ip1(n27325), .ip2(\LUT[110][4] ), .op(n25486) );
  nand4_1 U29495 ( .ip1(n25489), .ip2(n25488), .ip3(n25487), .ip4(n25486), 
        .op(n25490) );
  not_ab_or_c_or_d U29496 ( .ip1(\LUT[102][4] ), .ip2(n27326), .ip3(n25491), 
        .ip4(n25490), .op(n25495) );
  nand2_1 U29497 ( .ip1(n27370), .ip2(\LUT[100][4] ), .op(n25494) );
  nand2_1 U29498 ( .ip1(n27328), .ip2(\LUT[101][4] ), .op(n25493) );
  nand2_1 U29499 ( .ip1(n27327), .ip2(\LUT[103][4] ), .op(n25492) );
  nand4_1 U29500 ( .ip1(n25495), .ip2(n25494), .ip3(n25493), .ip4(n25492), 
        .op(n25496) );
  not_ab_or_c_or_d U29501 ( .ip1(\LUT[99][4] ), .ip2(n27156), .ip3(n25497), 
        .ip4(n25496), .op(n25498) );
  nor2_1 U29502 ( .ip1(n25498), .ip2(n27371), .op(n25511) );
  nand2_1 U29503 ( .ip1(n27582), .ip2(\LUT[115][4] ), .op(n25502) );
  nand2_1 U29504 ( .ip1(n27298), .ip2(\LUT[117][4] ), .op(n25501) );
  nand2_1 U29505 ( .ip1(n27299), .ip2(\LUT[118][4] ), .op(n25500) );
  nand2_1 U29506 ( .ip1(n27300), .ip2(\LUT[119][4] ), .op(n25499) );
  nand4_1 U29507 ( .ip1(n25502), .ip2(n25501), .ip3(n25500), .ip4(n25499), 
        .op(n25503) );
  or2_1 U29508 ( .ip1(n27297), .ip2(n25503), .op(n25505) );
  or2_1 U29509 ( .ip1(\LUT[116][4] ), .ip2(n25503), .op(n25504) );
  nand2_1 U29510 ( .ip1(n25505), .ip2(n25504), .op(n25509) );
  nand2_1 U29511 ( .ip1(n27165), .ip2(\LUT[108][4] ), .op(n25508) );
  nand2_1 U29512 ( .ip1(n27289), .ip2(\LUT[112][4] ), .op(n25507) );
  nand2_1 U29513 ( .ip1(n27305), .ip2(\LUT[114][4] ), .op(n25506) );
  nand4_1 U29514 ( .ip1(n25509), .ip2(n25508), .ip3(n25507), .ip4(n25506), 
        .op(n25510) );
  not_ab_or_c_or_d U29515 ( .ip1(n27583), .ip2(\LUT[113][4] ), .ip3(n25511), 
        .ip4(n25510), .op(n25629) );
  and2_1 U29516 ( .ip1(n27534), .ip2(\LUT[65][4] ), .op(n25517) );
  nand2_1 U29517 ( .ip1(n27548), .ip2(\LUT[67][4] ), .op(n25515) );
  nand2_1 U29518 ( .ip1(n27537), .ip2(\LUT[68][4] ), .op(n25514) );
  nand2_1 U29519 ( .ip1(n27535), .ip2(\LUT[69][4] ), .op(n25513) );
  nand2_1 U29520 ( .ip1(n27536), .ip2(\LUT[70][4] ), .op(n25512) );
  nand4_1 U29521 ( .ip1(n25515), .ip2(n25514), .ip3(n25513), .ip4(n25512), 
        .op(n25516) );
  not_ab_or_c_or_d U29522 ( .ip1(n27542), .ip2(\LUT[66][4] ), .ip3(n25517), 
        .ip4(n25516), .op(n25521) );
  nand2_1 U29523 ( .ip1(n27547), .ip2(\LUT[64][4] ), .op(n25520) );
  nand2_1 U29524 ( .ip1(n27546), .ip2(\LUT[59][4] ), .op(n25519) );
  nand2_1 U29525 ( .ip1(n27563), .ip2(\LUT[62][4] ), .op(n25518) );
  nand4_1 U29526 ( .ip1(n25521), .ip2(n25520), .ip3(n25519), .ip4(n25518), 
        .op(n25527) );
  nand2_1 U29527 ( .ip1(n27397), .ip2(\LUT[58][4] ), .op(n25525) );
  nand2_1 U29528 ( .ip1(n27555), .ip2(\LUT[61][4] ), .op(n25524) );
  nand2_1 U29529 ( .ip1(n27556), .ip2(\LUT[63][4] ), .op(n25523) );
  nand2_1 U29530 ( .ip1(n27554), .ip2(\LUT[60][4] ), .op(n25522) );
  nand4_1 U29531 ( .ip1(n25525), .ip2(n25524), .ip3(n25523), .ip4(n25522), 
        .op(n25526) );
  not_ab_or_c_or_d U29532 ( .ip1(n27553), .ip2(\LUT[57][4] ), .ip3(n25527), 
        .ip4(n25526), .op(n25528) );
  or2_1 U29533 ( .ip1(n25528), .ip2(n27265), .op(n25606) );
  nand2_1 U29534 ( .ip1(\LUT[27][4] ), .ip2(n27398), .op(n25531) );
  nand2_1 U29535 ( .ip1(n27400), .ip2(\LUT[28][4] ), .op(n25530) );
  nand2_1 U29536 ( .ip1(n27399), .ip2(\LUT[26][4] ), .op(n25529) );
  nand3_1 U29537 ( .ip1(n25531), .ip2(n25530), .ip3(n25529), .op(n25536) );
  nand2_1 U29538 ( .ip1(n27404), .ip2(\LUT[24][4] ), .op(n25534) );
  nand2_1 U29539 ( .ip1(n27405), .ip2(\LUT[25][4] ), .op(n25533) );
  nand2_1 U29540 ( .ip1(n27406), .ip2(\LUT[23][4] ), .op(n25532) );
  nand3_1 U29541 ( .ip1(n25534), .ip2(n25533), .ip3(n25532), .op(n25535) );
  not_ab_or_c_or_d U29542 ( .ip1(n27459), .ip2(\LUT[17][4] ), .ip3(n25536), 
        .ip4(n25535), .op(n25565) );
  nand2_1 U29543 ( .ip1(\LUT[2][4] ), .ip2(n27413), .op(n25538) );
  nand2_1 U29544 ( .ip1(\LUT[3][4] ), .ip2(n27414), .op(n25537) );
  nand2_1 U29545 ( .ip1(n25538), .ip2(n25537), .op(n25554) );
  nand2_1 U29546 ( .ip1(n27417), .ip2(\LUT[7][4] ), .op(n25542) );
  nand2_1 U29547 ( .ip1(n27418), .ip2(\LUT[9][4] ), .op(n25541) );
  nand2_1 U29548 ( .ip1(n27420), .ip2(\LUT[13][4] ), .op(n25540) );
  nand2_1 U29549 ( .ip1(n27419), .ip2(\LUT[14][4] ), .op(n25539) );
  nand4_1 U29550 ( .ip1(n25542), .ip2(n25541), .ip3(n25540), .ip4(n25539), 
        .op(n25548) );
  nand2_1 U29551 ( .ip1(n27425), .ip2(\LUT[10][4] ), .op(n25546) );
  nand2_1 U29552 ( .ip1(n27427), .ip2(\LUT[12][4] ), .op(n25545) );
  nand2_1 U29553 ( .ip1(n27428), .ip2(\LUT[6][4] ), .op(n25544) );
  nand2_1 U29554 ( .ip1(n27426), .ip2(\LUT[8][4] ), .op(n25543) );
  nand4_1 U29555 ( .ip1(n25546), .ip2(n25545), .ip3(n25544), .ip4(n25543), 
        .op(n25547) );
  not_ab_or_c_or_d U29556 ( .ip1(n27435), .ip2(\LUT[11][4] ), .ip3(n25548), 
        .ip4(n25547), .op(n25552) );
  nand2_1 U29557 ( .ip1(n27445), .ip2(\LUT[1][4] ), .op(n25551) );
  nand2_1 U29558 ( .ip1(n27438), .ip2(\LUT[5][4] ), .op(n25550) );
  nand2_1 U29559 ( .ip1(n27437), .ip2(\LUT[4][4] ), .op(n25549) );
  nand4_1 U29560 ( .ip1(n25552), .ip2(n25551), .ip3(n25550), .ip4(n25549), 
        .op(n25553) );
  not_ab_or_c_or_d U29561 ( .ip1(n27436), .ip2(\LUT[0][4] ), .ip3(n25554), 
        .ip4(n25553), .op(n25555) );
  nor2_1 U29562 ( .ip1(n25555), .ip2(n27446), .op(n25561) );
  nand2_1 U29563 ( .ip1(n27451), .ip2(\LUT[16][4] ), .op(n25559) );
  nand2_1 U29564 ( .ip1(n27449), .ip2(\LUT[20][4] ), .op(n25558) );
  nand2_1 U29565 ( .ip1(n27448), .ip2(\LUT[18][4] ), .op(n25557) );
  nand2_1 U29566 ( .ip1(n27450), .ip2(\LUT[21][4] ), .op(n25556) );
  nand4_1 U29567 ( .ip1(n25559), .ip2(n25558), .ip3(n25557), .ip4(n25556), 
        .op(n25560) );
  not_ab_or_c_or_d U29568 ( .ip1(\LUT[15][4] ), .ip2(n27458), .ip3(n25561), 
        .ip4(n25560), .op(n25564) );
  nand2_1 U29569 ( .ip1(n27460), .ip2(\LUT[19][4] ), .op(n25563) );
  nand2_1 U29570 ( .ip1(n27412), .ip2(\LUT[22][4] ), .op(n25562) );
  nand4_1 U29571 ( .ip1(n25565), .ip2(n25564), .ip3(n25563), .ip4(n25562), 
        .op(n25603) );
  nand2_1 U29572 ( .ip1(n27498), .ip2(\LUT[48][4] ), .op(n25569) );
  nand2_1 U29573 ( .ip1(n27499), .ip2(\LUT[49][4] ), .op(n25568) );
  nand2_1 U29574 ( .ip1(n27501), .ip2(\LUT[52][4] ), .op(n25567) );
  nand2_1 U29575 ( .ip1(n27500), .ip2(\LUT[53][4] ), .op(n25566) );
  nand4_1 U29576 ( .ip1(n25569), .ip2(n25568), .ip3(n25567), .ip4(n25566), 
        .op(n25581) );
  and2_1 U29577 ( .ip1(n27518), .ip2(\LUT[44][4] ), .op(n25575) );
  nand2_1 U29578 ( .ip1(n27508), .ip2(\LUT[55][4] ), .op(n25573) );
  nand2_1 U29579 ( .ip1(n27509), .ip2(\LUT[56][4] ), .op(n25572) );
  nand2_1 U29580 ( .ip1(n27507), .ip2(\LUT[54][4] ), .op(n25571) );
  nand2_1 U29581 ( .ip1(n27510), .ip2(\LUT[51][4] ), .op(n25570) );
  nand4_1 U29582 ( .ip1(n25573), .ip2(n25572), .ip3(n25571), .ip4(n25570), 
        .op(n25574) );
  not_ab_or_c_or_d U29583 ( .ip1(n27517), .ip2(\LUT[50][4] ), .ip3(n25575), 
        .ip4(n25574), .op(n25579) );
  nand2_1 U29584 ( .ip1(n27506), .ip2(\LUT[45][4] ), .op(n25578) );
  nand2_1 U29585 ( .ip1(n27519), .ip2(\LUT[43][4] ), .op(n25577) );
  nand2_1 U29586 ( .ip1(n27520), .ip2(\LUT[47][4] ), .op(n25576) );
  nand4_1 U29587 ( .ip1(n25579), .ip2(n25578), .ip3(n25577), .ip4(n25576), 
        .op(n25580) );
  not_ab_or_c_or_d U29588 ( .ip1(n27527), .ip2(\LUT[46][4] ), .ip3(n25581), 
        .ip4(n25580), .op(n25582) );
  nor2_1 U29589 ( .ip1(n25582), .ip2(n27528), .op(n25602) );
  nand2_1 U29590 ( .ip1(\LUT[31][4] ), .ip2(n27465), .op(n25584) );
  nand2_1 U29591 ( .ip1(\LUT[30][4] ), .ip2(n27466), .op(n25583) );
  nand2_1 U29592 ( .ip1(n25584), .ip2(n25583), .op(n25599) );
  nand2_1 U29593 ( .ip1(n27469), .ip2(\LUT[39][4] ), .op(n25588) );
  nand2_1 U29594 ( .ip1(n27470), .ip2(\LUT[38][4] ), .op(n25587) );
  nand2_1 U29595 ( .ip1(n27471), .ip2(\LUT[41][4] ), .op(n25586) );
  nand2_1 U29596 ( .ip1(n27472), .ip2(\LUT[42][4] ), .op(n25585) );
  nand4_1 U29597 ( .ip1(n25588), .ip2(n25587), .ip3(n25586), .ip4(n25585), 
        .op(n25593) );
  nand2_1 U29598 ( .ip1(\LUT[36][4] ), .ip2(n27477), .op(n25591) );
  nand2_1 U29599 ( .ip1(n27478), .ip2(\LUT[37][4] ), .op(n25590) );
  nand2_1 U29600 ( .ip1(n27488), .ip2(\LUT[33][4] ), .op(n25589) );
  nand3_1 U29601 ( .ip1(n25591), .ip2(n25590), .ip3(n25589), .op(n25592) );
  not_ab_or_c_or_d U29602 ( .ip1(n27485), .ip2(\LUT[40][4] ), .ip3(n25593), 
        .ip4(n25592), .op(n25597) );
  nand2_1 U29603 ( .ip1(n27486), .ip2(\LUT[34][4] ), .op(n25596) );
  nand2_1 U29604 ( .ip1(n27487), .ip2(\LUT[35][4] ), .op(n25595) );
  nand2_1 U29605 ( .ip1(n27479), .ip2(\LUT[32][4] ), .op(n25594) );
  nand4_1 U29606 ( .ip1(n25597), .ip2(n25596), .ip3(n25595), .ip4(n25594), 
        .op(n25598) );
  not_ab_or_c_or_d U29607 ( .ip1(n27495), .ip2(\LUT[29][4] ), .ip3(n25599), 
        .ip4(n25598), .op(n25600) );
  nor2_1 U29608 ( .ip1(n25600), .ip2(n27496), .op(n25601) );
  not_ab_or_c_or_d U29609 ( .ip1(n27533), .ip2(n25603), .ip3(n25602), .ip4(
        n25601), .op(n25604) );
  or2_1 U29610 ( .ip1(n25604), .ip2(n27265), .op(n25605) );
  nand2_1 U29611 ( .ip1(n25606), .ip2(n25605), .op(n25620) );
  nand2_1 U29612 ( .ip1(n27391), .ip2(\LUT[75][4] ), .op(n25618) );
  nand2_1 U29613 ( .ip1(n27373), .ip2(\LUT[82][4] ), .op(n25610) );
  nand2_1 U29614 ( .ip1(n27374), .ip2(\LUT[81][4] ), .op(n25609) );
  nand2_1 U29615 ( .ip1(n27375), .ip2(\LUT[84][4] ), .op(n25608) );
  nand2_1 U29616 ( .ip1(n27376), .ip2(\LUT[83][4] ), .op(n25607) );
  nand4_1 U29617 ( .ip1(n25610), .ip2(n25609), .ip3(n25608), .ip4(n25607), 
        .op(n25615) );
  nand2_1 U29618 ( .ip1(n27381), .ip2(\LUT[78][4] ), .op(n25613) );
  nand2_1 U29619 ( .ip1(n27382), .ip2(\LUT[79][4] ), .op(n25612) );
  nand2_1 U29620 ( .ip1(n27383), .ip2(\LUT[77][4] ), .op(n25611) );
  nand3_1 U29621 ( .ip1(n25613), .ip2(n25612), .ip3(n25611), .op(n25614) );
  not_ab_or_c_or_d U29622 ( .ip1(n27389), .ip2(\LUT[80][4] ), .ip3(n25615), 
        .ip4(n25614), .op(n25617) );
  nand2_1 U29623 ( .ip1(n27392), .ip2(\LUT[74][4] ), .op(n25616) );
  nand3_1 U29624 ( .ip1(n25618), .ip2(n25617), .ip3(n25616), .op(n25619) );
  not_ab_or_c_or_d U29625 ( .ip1(n27390), .ip2(\LUT[76][4] ), .ip3(n25620), 
        .ip4(n25619), .op(n25624) );
  nand2_1 U29626 ( .ip1(n27576), .ip2(\LUT[71][4] ), .op(n25623) );
  nand2_1 U29627 ( .ip1(n27570), .ip2(\LUT[72][4] ), .op(n25622) );
  nand2_1 U29628 ( .ip1(n27569), .ip2(\LUT[73][4] ), .op(n25621) );
  nand4_1 U29629 ( .ip1(n25624), .ip2(n25623), .ip3(n25622), .ip4(n25621), 
        .op(n25625) );
  nand2_1 U29630 ( .ip1(n27288), .ip2(n25625), .op(n25628) );
  nand2_1 U29631 ( .ip1(n27581), .ip2(\LUT[106][4] ), .op(n25627) );
  nand2_1 U29632 ( .ip1(n27172), .ip2(\LUT[111][4] ), .op(n25626) );
  nand4_1 U29633 ( .ip1(n25629), .ip2(n25628), .ip3(n25627), .ip4(n25626), 
        .op(n25630) );
  nand2_1 U29634 ( .ip1(n27589), .ip2(n25630), .op(n25632) );
  nand2_1 U29635 ( .ip1(sig_out[4]), .ip2(n27590), .op(n25631) );
  nand2_1 U29636 ( .ip1(n25632), .ip2(n25631), .op(n13461) );
  nand2_1 U29637 ( .ip1(n27333), .ip2(\LUT[95][5] ), .op(n25636) );
  nand2_1 U29638 ( .ip1(n27334), .ip2(\LUT[94][5] ), .op(n25635) );
  nand2_1 U29639 ( .ip1(n27336), .ip2(\LUT[97][5] ), .op(n25634) );
  nand2_1 U29640 ( .ip1(n27335), .ip2(\LUT[98][5] ), .op(n25633) );
  nand4_1 U29641 ( .ip1(n25636), .ip2(n25635), .ip3(n25634), .ip4(n25633), 
        .op(n25641) );
  nand2_1 U29642 ( .ip1(n27341), .ip2(\LUT[93][5] ), .op(n25639) );
  nand2_1 U29643 ( .ip1(n27342), .ip2(\LUT[92][5] ), .op(n25638) );
  nand2_1 U29644 ( .ip1(n27343), .ip2(\LUT[91][5] ), .op(n25637) );
  nand3_1 U29645 ( .ip1(n25639), .ip2(n25638), .ip3(n25637), .op(n25640) );
  not_ab_or_c_or_d U29646 ( .ip1(n27349), .ip2(\LUT[96][5] ), .ip3(n25641), 
        .ip4(n25640), .op(n25645) );
  nand2_1 U29647 ( .ip1(n27350), .ip2(\LUT[89][5] ), .op(n25644) );
  nand2_1 U29648 ( .ip1(n27351), .ip2(\LUT[90][5] ), .op(n25643) );
  nand2_1 U29649 ( .ip1(n27352), .ip2(\LUT[88][5] ), .op(n25642) );
  nand4_1 U29650 ( .ip1(n25645), .ip2(n25644), .ip3(n25643), .ip4(n25642), 
        .op(n25649) );
  nand2_1 U29651 ( .ip1(\LUT[85][5] ), .ip2(n27357), .op(n25647) );
  nand2_1 U29652 ( .ip1(\LUT[86][5] ), .ip2(n27358), .op(n25646) );
  nand2_1 U29653 ( .ip1(n25647), .ip2(n25646), .op(n25648) );
  not_ab_or_c_or_d U29654 ( .ip1(n27363), .ip2(\LUT[87][5] ), .ip3(n25649), 
        .ip4(n25648), .op(n25650) );
  nor2_1 U29655 ( .ip1(n25650), .ip2(n27142), .op(n25662) );
  and2_1 U29656 ( .ip1(n27317), .ip2(\LUT[105][5] ), .op(n25656) );
  nand2_1 U29657 ( .ip1(n27318), .ip2(\LUT[107][5] ), .op(n25654) );
  nand2_1 U29658 ( .ip1(n27319), .ip2(\LUT[104][5] ), .op(n25653) );
  nand2_1 U29659 ( .ip1(n27325), .ip2(\LUT[110][5] ), .op(n25652) );
  nand2_1 U29660 ( .ip1(n27309), .ip2(\LUT[109][5] ), .op(n25651) );
  nand4_1 U29661 ( .ip1(n25654), .ip2(n25653), .ip3(n25652), .ip4(n25651), 
        .op(n25655) );
  not_ab_or_c_or_d U29662 ( .ip1(\LUT[102][5] ), .ip2(n27326), .ip3(n25656), 
        .ip4(n25655), .op(n25660) );
  nand2_1 U29663 ( .ip1(n27370), .ip2(\LUT[100][5] ), .op(n25659) );
  nand2_1 U29664 ( .ip1(n27328), .ip2(\LUT[101][5] ), .op(n25658) );
  nand2_1 U29665 ( .ip1(n27327), .ip2(\LUT[103][5] ), .op(n25657) );
  nand4_1 U29666 ( .ip1(n25660), .ip2(n25659), .ip3(n25658), .ip4(n25657), 
        .op(n25661) );
  not_ab_or_c_or_d U29667 ( .ip1(\LUT[99][5] ), .ip2(n27156), .ip3(n25662), 
        .ip4(n25661), .op(n25663) );
  nor2_1 U29668 ( .ip1(n25663), .ip2(n27371), .op(n25676) );
  nand2_1 U29669 ( .ip1(n27582), .ip2(\LUT[115][5] ), .op(n25667) );
  nand2_1 U29670 ( .ip1(n27298), .ip2(\LUT[117][5] ), .op(n25666) );
  nand2_1 U29671 ( .ip1(n27299), .ip2(\LUT[118][5] ), .op(n25665) );
  nand2_1 U29672 ( .ip1(n27300), .ip2(\LUT[119][5] ), .op(n25664) );
  nand4_1 U29673 ( .ip1(n25667), .ip2(n25666), .ip3(n25665), .ip4(n25664), 
        .op(n25668) );
  or2_1 U29674 ( .ip1(n27297), .ip2(n25668), .op(n25670) );
  or2_1 U29675 ( .ip1(\LUT[116][5] ), .ip2(n25668), .op(n25669) );
  nand2_1 U29676 ( .ip1(n25670), .ip2(n25669), .op(n25674) );
  nand2_1 U29677 ( .ip1(n27289), .ip2(\LUT[112][5] ), .op(n25673) );
  nand2_1 U29678 ( .ip1(n27165), .ip2(\LUT[108][5] ), .op(n25672) );
  nand2_1 U29679 ( .ip1(n27305), .ip2(\LUT[114][5] ), .op(n25671) );
  nand4_1 U29680 ( .ip1(n25674), .ip2(n25673), .ip3(n25672), .ip4(n25671), 
        .op(n25675) );
  not_ab_or_c_or_d U29681 ( .ip1(n27583), .ip2(\LUT[113][5] ), .ip3(n25676), 
        .ip4(n25675), .op(n25794) );
  and2_1 U29682 ( .ip1(n27548), .ip2(\LUT[67][5] ), .op(n25682) );
  nand2_1 U29683 ( .ip1(n27534), .ip2(\LUT[65][5] ), .op(n25680) );
  nand2_1 U29684 ( .ip1(n27535), .ip2(\LUT[69][5] ), .op(n25679) );
  nand2_1 U29685 ( .ip1(n27536), .ip2(\LUT[70][5] ), .op(n25678) );
  nand2_1 U29686 ( .ip1(n27537), .ip2(\LUT[68][5] ), .op(n25677) );
  nand4_1 U29687 ( .ip1(n25680), .ip2(n25679), .ip3(n25678), .ip4(n25677), 
        .op(n25681) );
  not_ab_or_c_or_d U29688 ( .ip1(n27542), .ip2(\LUT[66][5] ), .ip3(n25682), 
        .ip4(n25681), .op(n25686) );
  nand2_1 U29689 ( .ip1(n27546), .ip2(\LUT[59][5] ), .op(n25685) );
  nand2_1 U29690 ( .ip1(n27547), .ip2(\LUT[64][5] ), .op(n25684) );
  nand2_1 U29691 ( .ip1(n27555), .ip2(\LUT[61][5] ), .op(n25683) );
  nand4_1 U29692 ( .ip1(n25686), .ip2(n25685), .ip3(n25684), .ip4(n25683), 
        .op(n25692) );
  nand2_1 U29693 ( .ip1(n27553), .ip2(\LUT[57][5] ), .op(n25690) );
  nand2_1 U29694 ( .ip1(n27563), .ip2(\LUT[62][5] ), .op(n25689) );
  nand2_1 U29695 ( .ip1(n27556), .ip2(\LUT[63][5] ), .op(n25688) );
  nand2_1 U29696 ( .ip1(n27554), .ip2(\LUT[60][5] ), .op(n25687) );
  nand4_1 U29697 ( .ip1(n25690), .ip2(n25689), .ip3(n25688), .ip4(n25687), 
        .op(n25691) );
  not_ab_or_c_or_d U29698 ( .ip1(n27397), .ip2(\LUT[58][5] ), .ip3(n25692), 
        .ip4(n25691), .op(n25693) );
  or2_1 U29699 ( .ip1(n25693), .ip2(n27265), .op(n25771) );
  nand2_1 U29700 ( .ip1(\LUT[27][5] ), .ip2(n27398), .op(n25696) );
  nand2_1 U29701 ( .ip1(n27399), .ip2(\LUT[26][5] ), .op(n25695) );
  nand2_1 U29702 ( .ip1(n27400), .ip2(\LUT[28][5] ), .op(n25694) );
  nand3_1 U29703 ( .ip1(n25696), .ip2(n25695), .ip3(n25694), .op(n25701) );
  nand2_1 U29704 ( .ip1(\LUT[24][5] ), .ip2(n27404), .op(n25699) );
  nand2_1 U29705 ( .ip1(n27405), .ip2(\LUT[25][5] ), .op(n25698) );
  nand2_1 U29706 ( .ip1(n27406), .ip2(\LUT[23][5] ), .op(n25697) );
  nand3_1 U29707 ( .ip1(n25699), .ip2(n25698), .ip3(n25697), .op(n25700) );
  not_ab_or_c_or_d U29708 ( .ip1(n27459), .ip2(\LUT[17][5] ), .ip3(n25701), 
        .ip4(n25700), .op(n25730) );
  nand2_1 U29709 ( .ip1(\LUT[2][5] ), .ip2(n27413), .op(n25703) );
  nand2_1 U29710 ( .ip1(\LUT[3][5] ), .ip2(n27414), .op(n25702) );
  nand2_1 U29711 ( .ip1(n25703), .ip2(n25702), .op(n25719) );
  nand2_1 U29712 ( .ip1(n27428), .ip2(\LUT[6][5] ), .op(n25707) );
  nand2_1 U29713 ( .ip1(n27427), .ip2(\LUT[12][5] ), .op(n25706) );
  nand2_1 U29714 ( .ip1(n27420), .ip2(\LUT[13][5] ), .op(n25705) );
  nand2_1 U29715 ( .ip1(n27419), .ip2(\LUT[14][5] ), .op(n25704) );
  nand4_1 U29716 ( .ip1(n25707), .ip2(n25706), .ip3(n25705), .ip4(n25704), 
        .op(n25713) );
  nand2_1 U29717 ( .ip1(n27426), .ip2(\LUT[8][5] ), .op(n25711) );
  nand2_1 U29718 ( .ip1(n27417), .ip2(\LUT[7][5] ), .op(n25710) );
  nand2_1 U29719 ( .ip1(n27425), .ip2(\LUT[10][5] ), .op(n25709) );
  nand2_1 U29720 ( .ip1(n27435), .ip2(\LUT[11][5] ), .op(n25708) );
  nand4_1 U29721 ( .ip1(n25711), .ip2(n25710), .ip3(n25709), .ip4(n25708), 
        .op(n25712) );
  not_ab_or_c_or_d U29722 ( .ip1(n27418), .ip2(\LUT[9][5] ), .ip3(n25713), 
        .ip4(n25712), .op(n25717) );
  nand2_1 U29723 ( .ip1(n27445), .ip2(\LUT[1][5] ), .op(n25716) );
  nand2_1 U29724 ( .ip1(n27438), .ip2(\LUT[5][5] ), .op(n25715) );
  nand2_1 U29725 ( .ip1(n27437), .ip2(\LUT[4][5] ), .op(n25714) );
  nand4_1 U29726 ( .ip1(n25717), .ip2(n25716), .ip3(n25715), .ip4(n25714), 
        .op(n25718) );
  not_ab_or_c_or_d U29727 ( .ip1(n27436), .ip2(\LUT[0][5] ), .ip3(n25719), 
        .ip4(n25718), .op(n25720) );
  nor2_1 U29728 ( .ip1(n25720), .ip2(n27446), .op(n25726) );
  nand2_1 U29729 ( .ip1(n27449), .ip2(\LUT[20][5] ), .op(n25724) );
  nand2_1 U29730 ( .ip1(n27450), .ip2(\LUT[21][5] ), .op(n25723) );
  nand2_1 U29731 ( .ip1(n27448), .ip2(\LUT[18][5] ), .op(n25722) );
  nand2_1 U29732 ( .ip1(n27451), .ip2(\LUT[16][5] ), .op(n25721) );
  nand4_1 U29733 ( .ip1(n25724), .ip2(n25723), .ip3(n25722), .ip4(n25721), 
        .op(n25725) );
  not_ab_or_c_or_d U29734 ( .ip1(\LUT[15][5] ), .ip2(n27458), .ip3(n25726), 
        .ip4(n25725), .op(n25729) );
  nand2_1 U29735 ( .ip1(n27412), .ip2(\LUT[22][5] ), .op(n25728) );
  nand2_1 U29736 ( .ip1(n27460), .ip2(\LUT[19][5] ), .op(n25727) );
  nand4_1 U29737 ( .ip1(n25730), .ip2(n25729), .ip3(n25728), .ip4(n25727), 
        .op(n25768) );
  nand2_1 U29738 ( .ip1(\LUT[31][5] ), .ip2(n27465), .op(n25732) );
  nand2_1 U29739 ( .ip1(\LUT[30][5] ), .ip2(n27466), .op(n25731) );
  nand2_1 U29740 ( .ip1(n25732), .ip2(n25731), .op(n25747) );
  nand2_1 U29741 ( .ip1(n27470), .ip2(\LUT[38][5] ), .op(n25736) );
  nand2_1 U29742 ( .ip1(n27469), .ip2(\LUT[39][5] ), .op(n25735) );
  nand2_1 U29743 ( .ip1(n27471), .ip2(\LUT[41][5] ), .op(n25734) );
  nand2_1 U29744 ( .ip1(n27472), .ip2(\LUT[42][5] ), .op(n25733) );
  nand4_1 U29745 ( .ip1(n25736), .ip2(n25735), .ip3(n25734), .ip4(n25733), 
        .op(n25741) );
  nand2_1 U29746 ( .ip1(n27477), .ip2(\LUT[36][5] ), .op(n25739) );
  nand2_1 U29747 ( .ip1(n27478), .ip2(\LUT[37][5] ), .op(n25738) );
  nand2_1 U29748 ( .ip1(n27479), .ip2(\LUT[32][5] ), .op(n25737) );
  nand3_1 U29749 ( .ip1(n25739), .ip2(n25738), .ip3(n25737), .op(n25740) );
  not_ab_or_c_or_d U29750 ( .ip1(n27485), .ip2(\LUT[40][5] ), .ip3(n25741), 
        .ip4(n25740), .op(n25745) );
  nand2_1 U29751 ( .ip1(n27487), .ip2(\LUT[35][5] ), .op(n25744) );
  nand2_1 U29752 ( .ip1(n27486), .ip2(\LUT[34][5] ), .op(n25743) );
  nand2_1 U29753 ( .ip1(n27488), .ip2(\LUT[33][5] ), .op(n25742) );
  nand4_1 U29754 ( .ip1(n25745), .ip2(n25744), .ip3(n25743), .ip4(n25742), 
        .op(n25746) );
  not_ab_or_c_or_d U29755 ( .ip1(n27495), .ip2(\LUT[29][5] ), .ip3(n25747), 
        .ip4(n25746), .op(n25748) );
  nor2_1 U29756 ( .ip1(n25748), .ip2(n27496), .op(n25767) );
  nand2_1 U29757 ( .ip1(n27499), .ip2(\LUT[49][5] ), .op(n25752) );
  nand2_1 U29758 ( .ip1(n27498), .ip2(\LUT[48][5] ), .op(n25751) );
  nand2_1 U29759 ( .ip1(n27500), .ip2(\LUT[53][5] ), .op(n25750) );
  nand2_1 U29760 ( .ip1(n27501), .ip2(\LUT[52][5] ), .op(n25749) );
  nand4_1 U29761 ( .ip1(n25752), .ip2(n25751), .ip3(n25750), .ip4(n25749), 
        .op(n25764) );
  and2_1 U29762 ( .ip1(n27506), .ip2(\LUT[45][5] ), .op(n25758) );
  nand2_1 U29763 ( .ip1(n27507), .ip2(\LUT[54][5] ), .op(n25756) );
  nand2_1 U29764 ( .ip1(n27509), .ip2(\LUT[56][5] ), .op(n25755) );
  nand2_1 U29765 ( .ip1(n27508), .ip2(\LUT[55][5] ), .op(n25754) );
  nand2_1 U29766 ( .ip1(n27510), .ip2(\LUT[51][5] ), .op(n25753) );
  nand4_1 U29767 ( .ip1(n25756), .ip2(n25755), .ip3(n25754), .ip4(n25753), 
        .op(n25757) );
  not_ab_or_c_or_d U29768 ( .ip1(n27517), .ip2(\LUT[50][5] ), .ip3(n25758), 
        .ip4(n25757), .op(n25762) );
  nand2_1 U29769 ( .ip1(n27518), .ip2(\LUT[44][5] ), .op(n25761) );
  nand2_1 U29770 ( .ip1(n27519), .ip2(\LUT[43][5] ), .op(n25760) );
  nand2_1 U29771 ( .ip1(n27520), .ip2(\LUT[47][5] ), .op(n25759) );
  nand4_1 U29772 ( .ip1(n25762), .ip2(n25761), .ip3(n25760), .ip4(n25759), 
        .op(n25763) );
  not_ab_or_c_or_d U29773 ( .ip1(n27527), .ip2(\LUT[46][5] ), .ip3(n25764), 
        .ip4(n25763), .op(n25765) );
  nor2_1 U29774 ( .ip1(n25765), .ip2(n27528), .op(n25766) );
  not_ab_or_c_or_d U29775 ( .ip1(n27533), .ip2(n25768), .ip3(n25767), .ip4(
        n25766), .op(n25769) );
  or2_1 U29776 ( .ip1(n25769), .ip2(n27265), .op(n25770) );
  nand2_1 U29777 ( .ip1(n25771), .ip2(n25770), .op(n25785) );
  nand2_1 U29778 ( .ip1(n27391), .ip2(\LUT[75][5] ), .op(n25783) );
  nand2_1 U29779 ( .ip1(n27373), .ip2(\LUT[82][5] ), .op(n25775) );
  nand2_1 U29780 ( .ip1(n27374), .ip2(\LUT[81][5] ), .op(n25774) );
  nand2_1 U29781 ( .ip1(n27375), .ip2(\LUT[84][5] ), .op(n25773) );
  nand2_1 U29782 ( .ip1(n27376), .ip2(\LUT[83][5] ), .op(n25772) );
  nand4_1 U29783 ( .ip1(n25775), .ip2(n25774), .ip3(n25773), .ip4(n25772), 
        .op(n25780) );
  nand2_1 U29784 ( .ip1(\LUT[78][5] ), .ip2(n27381), .op(n25778) );
  nand2_1 U29785 ( .ip1(n27382), .ip2(\LUT[79][5] ), .op(n25777) );
  nand2_1 U29786 ( .ip1(n27383), .ip2(\LUT[77][5] ), .op(n25776) );
  nand3_1 U29787 ( .ip1(n25778), .ip2(n25777), .ip3(n25776), .op(n25779) );
  not_ab_or_c_or_d U29788 ( .ip1(n27389), .ip2(\LUT[80][5] ), .ip3(n25780), 
        .ip4(n25779), .op(n25782) );
  nand2_1 U29789 ( .ip1(n27392), .ip2(\LUT[74][5] ), .op(n25781) );
  nand3_1 U29790 ( .ip1(n25783), .ip2(n25782), .ip3(n25781), .op(n25784) );
  not_ab_or_c_or_d U29791 ( .ip1(n27390), .ip2(\LUT[76][5] ), .ip3(n25785), 
        .ip4(n25784), .op(n25789) );
  nand2_1 U29792 ( .ip1(n27576), .ip2(\LUT[71][5] ), .op(n25788) );
  nand2_1 U29793 ( .ip1(n27570), .ip2(\LUT[72][5] ), .op(n25787) );
  nand2_1 U29794 ( .ip1(n27569), .ip2(\LUT[73][5] ), .op(n25786) );
  nand4_1 U29795 ( .ip1(n25789), .ip2(n25788), .ip3(n25787), .ip4(n25786), 
        .op(n25790) );
  nand2_1 U29796 ( .ip1(n27288), .ip2(n25790), .op(n25793) );
  nand2_1 U29797 ( .ip1(n27581), .ip2(\LUT[106][5] ), .op(n25792) );
  nand2_1 U29798 ( .ip1(n27172), .ip2(\LUT[111][5] ), .op(n25791) );
  nand4_1 U29799 ( .ip1(n25794), .ip2(n25793), .ip3(n25792), .ip4(n25791), 
        .op(n25795) );
  nand2_1 U29800 ( .ip1(n27589), .ip2(n25795), .op(n25797) );
  nand2_1 U29801 ( .ip1(sig_out[5]), .ip2(n27590), .op(n25796) );
  nand2_1 U29802 ( .ip1(n25797), .ip2(n25796), .op(n13460) );
  nand2_1 U29803 ( .ip1(n27333), .ip2(\LUT[95][6] ), .op(n25801) );
  nand2_1 U29804 ( .ip1(n27334), .ip2(\LUT[94][6] ), .op(n25800) );
  nand2_1 U29805 ( .ip1(n27336), .ip2(\LUT[97][6] ), .op(n25799) );
  nand2_1 U29806 ( .ip1(n27335), .ip2(\LUT[98][6] ), .op(n25798) );
  nand4_1 U29807 ( .ip1(n25801), .ip2(n25800), .ip3(n25799), .ip4(n25798), 
        .op(n25806) );
  nand2_1 U29808 ( .ip1(n27341), .ip2(\LUT[93][6] ), .op(n25804) );
  nand2_1 U29809 ( .ip1(n27342), .ip2(\LUT[92][6] ), .op(n25803) );
  nand2_1 U29810 ( .ip1(n27343), .ip2(\LUT[91][6] ), .op(n25802) );
  nand3_1 U29811 ( .ip1(n25804), .ip2(n25803), .ip3(n25802), .op(n25805) );
  not_ab_or_c_or_d U29812 ( .ip1(n27349), .ip2(\LUT[96][6] ), .ip3(n25806), 
        .ip4(n25805), .op(n25810) );
  nand2_1 U29813 ( .ip1(n27350), .ip2(\LUT[89][6] ), .op(n25809) );
  nand2_1 U29814 ( .ip1(n27351), .ip2(\LUT[90][6] ), .op(n25808) );
  nand2_1 U29815 ( .ip1(n27352), .ip2(\LUT[88][6] ), .op(n25807) );
  nand4_1 U29816 ( .ip1(n25810), .ip2(n25809), .ip3(n25808), .ip4(n25807), 
        .op(n25814) );
  nand2_1 U29817 ( .ip1(\LUT[85][6] ), .ip2(n27357), .op(n25812) );
  nand2_1 U29818 ( .ip1(\LUT[86][6] ), .ip2(n27358), .op(n25811) );
  nand2_1 U29819 ( .ip1(n25812), .ip2(n25811), .op(n25813) );
  not_ab_or_c_or_d U29820 ( .ip1(n27363), .ip2(\LUT[87][6] ), .ip3(n25814), 
        .ip4(n25813), .op(n25815) );
  nor2_1 U29821 ( .ip1(n25815), .ip2(n27142), .op(n25827) );
  and2_1 U29822 ( .ip1(n27317), .ip2(\LUT[105][6] ), .op(n25821) );
  nand2_1 U29823 ( .ip1(n27318), .ip2(\LUT[107][6] ), .op(n25819) );
  nand2_1 U29824 ( .ip1(n27319), .ip2(\LUT[104][6] ), .op(n25818) );
  nand2_1 U29825 ( .ip1(n27325), .ip2(\LUT[110][6] ), .op(n25817) );
  nand2_1 U29826 ( .ip1(n27309), .ip2(\LUT[109][6] ), .op(n25816) );
  nand4_1 U29827 ( .ip1(n25819), .ip2(n25818), .ip3(n25817), .ip4(n25816), 
        .op(n25820) );
  not_ab_or_c_or_d U29828 ( .ip1(\LUT[102][6] ), .ip2(n27326), .ip3(n25821), 
        .ip4(n25820), .op(n25825) );
  nand2_1 U29829 ( .ip1(n27370), .ip2(\LUT[100][6] ), .op(n25824) );
  nand2_1 U29830 ( .ip1(n27328), .ip2(\LUT[101][6] ), .op(n25823) );
  nand2_1 U29831 ( .ip1(n27327), .ip2(\LUT[103][6] ), .op(n25822) );
  nand4_1 U29832 ( .ip1(n25825), .ip2(n25824), .ip3(n25823), .ip4(n25822), 
        .op(n25826) );
  not_ab_or_c_or_d U29833 ( .ip1(\LUT[99][6] ), .ip2(n27156), .ip3(n25827), 
        .ip4(n25826), .op(n25828) );
  nor2_1 U29834 ( .ip1(n25828), .ip2(n27371), .op(n25841) );
  nand2_1 U29835 ( .ip1(n27582), .ip2(\LUT[115][6] ), .op(n25832) );
  nand2_1 U29836 ( .ip1(n27298), .ip2(\LUT[117][6] ), .op(n25831) );
  nand2_1 U29837 ( .ip1(n27299), .ip2(\LUT[118][6] ), .op(n25830) );
  nand2_1 U29838 ( .ip1(n27300), .ip2(\LUT[119][6] ), .op(n25829) );
  nand4_1 U29839 ( .ip1(n25832), .ip2(n25831), .ip3(n25830), .ip4(n25829), 
        .op(n25833) );
  or2_1 U29840 ( .ip1(n27297), .ip2(n25833), .op(n25835) );
  or2_1 U29841 ( .ip1(\LUT[116][6] ), .ip2(n25833), .op(n25834) );
  nand2_1 U29842 ( .ip1(n25835), .ip2(n25834), .op(n25839) );
  nand2_1 U29843 ( .ip1(n27289), .ip2(\LUT[112][6] ), .op(n25838) );
  nand2_1 U29844 ( .ip1(n27165), .ip2(\LUT[108][6] ), .op(n25837) );
  nand2_1 U29845 ( .ip1(n27305), .ip2(\LUT[114][6] ), .op(n25836) );
  nand4_1 U29846 ( .ip1(n25839), .ip2(n25838), .ip3(n25837), .ip4(n25836), 
        .op(n25840) );
  not_ab_or_c_or_d U29847 ( .ip1(n27583), .ip2(\LUT[113][6] ), .ip3(n25841), 
        .ip4(n25840), .op(n25961) );
  nand2_1 U29848 ( .ip1(n27373), .ip2(\LUT[82][6] ), .op(n25845) );
  nand2_1 U29849 ( .ip1(n27374), .ip2(\LUT[81][6] ), .op(n25844) );
  nand2_1 U29850 ( .ip1(n27375), .ip2(\LUT[84][6] ), .op(n25843) );
  nand2_1 U29851 ( .ip1(n27376), .ip2(\LUT[83][6] ), .op(n25842) );
  nand4_1 U29852 ( .ip1(n25845), .ip2(n25844), .ip3(n25843), .ip4(n25842), 
        .op(n25850) );
  nand2_1 U29853 ( .ip1(n27381), .ip2(\LUT[78][6] ), .op(n25848) );
  nand2_1 U29854 ( .ip1(n27382), .ip2(\LUT[79][6] ), .op(n25847) );
  nand2_1 U29855 ( .ip1(n27383), .ip2(\LUT[77][6] ), .op(n25846) );
  nand3_1 U29856 ( .ip1(n25848), .ip2(n25847), .ip3(n25846), .op(n25849) );
  not_ab_or_c_or_d U29857 ( .ip1(n27389), .ip2(\LUT[80][6] ), .ip3(n25850), 
        .ip4(n25849), .op(n25854) );
  nand2_1 U29858 ( .ip1(n27390), .ip2(\LUT[76][6] ), .op(n25853) );
  nand2_1 U29859 ( .ip1(n27391), .ip2(\LUT[75][6] ), .op(n25852) );
  nand2_1 U29860 ( .ip1(n27392), .ip2(\LUT[74][6] ), .op(n25851) );
  nand4_1 U29861 ( .ip1(n25854), .ip2(n25853), .ip3(n25852), .ip4(n25851), 
        .op(n25956) );
  nand2_1 U29862 ( .ip1(n27548), .ip2(\LUT[67][6] ), .op(n25858) );
  nand2_1 U29863 ( .ip1(n27537), .ip2(\LUT[68][6] ), .op(n25857) );
  nand2_1 U29864 ( .ip1(n27535), .ip2(\LUT[69][6] ), .op(n25856) );
  nand2_1 U29865 ( .ip1(n27536), .ip2(\LUT[70][6] ), .op(n25855) );
  nand4_1 U29866 ( .ip1(n25858), .ip2(n25857), .ip3(n25856), .ip4(n25855), 
        .op(n25863) );
  nand2_1 U29867 ( .ip1(n27547), .ip2(\LUT[64][6] ), .op(n25861) );
  nand2_1 U29868 ( .ip1(n27542), .ip2(\LUT[66][6] ), .op(n25860) );
  nand2_1 U29869 ( .ip1(n27534), .ip2(\LUT[65][6] ), .op(n25859) );
  nand3_1 U29870 ( .ip1(n25861), .ip2(n25860), .ip3(n25859), .op(n25862) );
  not_ab_or_c_or_d U29871 ( .ip1(n27556), .ip2(\LUT[63][6] ), .ip3(n25863), 
        .ip4(n25862), .op(n25950) );
  nand2_1 U29872 ( .ip1(\LUT[27][6] ), .ip2(n27398), .op(n25866) );
  nand2_1 U29873 ( .ip1(n27399), .ip2(\LUT[26][6] ), .op(n25865) );
  nand2_1 U29874 ( .ip1(n27400), .ip2(\LUT[28][6] ), .op(n25864) );
  nand3_1 U29875 ( .ip1(n25866), .ip2(n25865), .ip3(n25864), .op(n25871) );
  nand2_1 U29876 ( .ip1(n27404), .ip2(\LUT[24][6] ), .op(n25869) );
  nand2_1 U29877 ( .ip1(n27405), .ip2(\LUT[25][6] ), .op(n25868) );
  nand2_1 U29878 ( .ip1(n27406), .ip2(\LUT[23][6] ), .op(n25867) );
  nand3_1 U29879 ( .ip1(n25869), .ip2(n25868), .ip3(n25867), .op(n25870) );
  not_ab_or_c_or_d U29880 ( .ip1(n27459), .ip2(\LUT[17][6] ), .ip3(n25871), 
        .ip4(n25870), .op(n25900) );
  nand2_1 U29881 ( .ip1(\LUT[2][6] ), .ip2(n27413), .op(n25873) );
  nand2_1 U29882 ( .ip1(\LUT[3][6] ), .ip2(n27414), .op(n25872) );
  nand2_1 U29883 ( .ip1(n25873), .ip2(n25872), .op(n25889) );
  nand2_1 U29884 ( .ip1(n27418), .ip2(\LUT[9][6] ), .op(n25877) );
  nand2_1 U29885 ( .ip1(n27417), .ip2(\LUT[7][6] ), .op(n25876) );
  nand2_1 U29886 ( .ip1(n27420), .ip2(\LUT[13][6] ), .op(n25875) );
  nand2_1 U29887 ( .ip1(n27419), .ip2(\LUT[14][6] ), .op(n25874) );
  nand4_1 U29888 ( .ip1(n25877), .ip2(n25876), .ip3(n25875), .ip4(n25874), 
        .op(n25883) );
  nand2_1 U29889 ( .ip1(n27425), .ip2(\LUT[10][6] ), .op(n25881) );
  nand2_1 U29890 ( .ip1(n27427), .ip2(\LUT[12][6] ), .op(n25880) );
  nand2_1 U29891 ( .ip1(n27426), .ip2(\LUT[8][6] ), .op(n25879) );
  nand2_1 U29892 ( .ip1(n27428), .ip2(\LUT[6][6] ), .op(n25878) );
  nand4_1 U29893 ( .ip1(n25881), .ip2(n25880), .ip3(n25879), .ip4(n25878), 
        .op(n25882) );
  not_ab_or_c_or_d U29894 ( .ip1(n27435), .ip2(\LUT[11][6] ), .ip3(n25883), 
        .ip4(n25882), .op(n25887) );
  nand2_1 U29895 ( .ip1(n27445), .ip2(\LUT[1][6] ), .op(n25886) );
  nand2_1 U29896 ( .ip1(n27437), .ip2(\LUT[4][6] ), .op(n25885) );
  nand2_1 U29897 ( .ip1(n27438), .ip2(\LUT[5][6] ), .op(n25884) );
  nand4_1 U29898 ( .ip1(n25887), .ip2(n25886), .ip3(n25885), .ip4(n25884), 
        .op(n25888) );
  not_ab_or_c_or_d U29899 ( .ip1(n27436), .ip2(\LUT[0][6] ), .ip3(n25889), 
        .ip4(n25888), .op(n25890) );
  nor2_1 U29900 ( .ip1(n25890), .ip2(n27446), .op(n25896) );
  nand2_1 U29901 ( .ip1(n27451), .ip2(\LUT[16][6] ), .op(n25894) );
  nand2_1 U29902 ( .ip1(n27449), .ip2(\LUT[20][6] ), .op(n25893) );
  nand2_1 U29903 ( .ip1(n27448), .ip2(\LUT[18][6] ), .op(n25892) );
  nand2_1 U29904 ( .ip1(n27450), .ip2(\LUT[21][6] ), .op(n25891) );
  nand4_1 U29905 ( .ip1(n25894), .ip2(n25893), .ip3(n25892), .ip4(n25891), 
        .op(n25895) );
  not_ab_or_c_or_d U29906 ( .ip1(\LUT[15][6] ), .ip2(n27458), .ip3(n25896), 
        .ip4(n25895), .op(n25899) );
  nand2_1 U29907 ( .ip1(n27460), .ip2(\LUT[19][6] ), .op(n25898) );
  nand2_1 U29908 ( .ip1(n27412), .ip2(\LUT[22][6] ), .op(n25897) );
  nand4_1 U29909 ( .ip1(n25900), .ip2(n25899), .ip3(n25898), .ip4(n25897), 
        .op(n25946) );
  nand2_1 U29910 ( .ip1(n27486), .ip2(\LUT[34][6] ), .op(n25903) );
  nand2_1 U29911 ( .ip1(n27487), .ip2(\LUT[35][6] ), .op(n25902) );
  nand2_1 U29912 ( .ip1(n27488), .ip2(\LUT[33][6] ), .op(n25901) );
  nand3_1 U29913 ( .ip1(n25903), .ip2(n25902), .ip3(n25901), .op(n25917) );
  nand2_1 U29914 ( .ip1(n27466), .ip2(\LUT[30][6] ), .op(n25915) );
  nand2_1 U29915 ( .ip1(n27469), .ip2(\LUT[39][6] ), .op(n25907) );
  nand2_1 U29916 ( .ip1(n27470), .ip2(\LUT[38][6] ), .op(n25906) );
  nand2_1 U29917 ( .ip1(n27471), .ip2(\LUT[41][6] ), .op(n25905) );
  nand2_1 U29918 ( .ip1(n27472), .ip2(\LUT[42][6] ), .op(n25904) );
  nand4_1 U29919 ( .ip1(n25907), .ip2(n25906), .ip3(n25905), .ip4(n25904), 
        .op(n25912) );
  nand2_1 U29920 ( .ip1(n27477), .ip2(\LUT[36][6] ), .op(n25910) );
  nand2_1 U29921 ( .ip1(n27478), .ip2(\LUT[37][6] ), .op(n25909) );
  nand2_1 U29922 ( .ip1(n27479), .ip2(\LUT[32][6] ), .op(n25908) );
  nand3_1 U29923 ( .ip1(n25910), .ip2(n25909), .ip3(n25908), .op(n25911) );
  not_ab_or_c_or_d U29924 ( .ip1(n27485), .ip2(\LUT[40][6] ), .ip3(n25912), 
        .ip4(n25911), .op(n25914) );
  nand2_1 U29925 ( .ip1(n27465), .ip2(\LUT[31][6] ), .op(n25913) );
  nand3_1 U29926 ( .ip1(n25915), .ip2(n25914), .ip3(n25913), .op(n25916) );
  not_ab_or_c_or_d U29927 ( .ip1(n27495), .ip2(\LUT[29][6] ), .ip3(n25917), 
        .ip4(n25916), .op(n25919) );
  inv_1 U29928 ( .ip(n25918), .op(n26743) );
  nor2_1 U29929 ( .ip1(n25919), .ip2(n26743), .op(n25938) );
  nand2_1 U29930 ( .ip1(n27500), .ip2(\LUT[53][6] ), .op(n25923) );
  nand2_1 U29931 ( .ip1(n27510), .ip2(\LUT[51][6] ), .op(n25922) );
  nand2_1 U29932 ( .ip1(n27508), .ip2(\LUT[55][6] ), .op(n25921) );
  nand2_1 U29933 ( .ip1(n27509), .ip2(\LUT[56][6] ), .op(n25920) );
  nand4_1 U29934 ( .ip1(n25923), .ip2(n25922), .ip3(n25921), .ip4(n25920), 
        .op(n25924) );
  or2_1 U29935 ( .ip1(n27520), .ip2(n25924), .op(n25926) );
  or2_1 U29936 ( .ip1(\LUT[47][6] ), .ip2(n25924), .op(n25925) );
  nand2_1 U29937 ( .ip1(n25926), .ip2(n25925), .op(n25936) );
  and2_1 U29938 ( .ip1(n27518), .ip2(\LUT[44][6] ), .op(n25932) );
  nand2_1 U29939 ( .ip1(n27498), .ip2(\LUT[48][6] ), .op(n25930) );
  nand2_1 U29940 ( .ip1(n27499), .ip2(\LUT[49][6] ), .op(n25929) );
  nand2_1 U29941 ( .ip1(n27507), .ip2(\LUT[54][6] ), .op(n25928) );
  nand2_1 U29942 ( .ip1(n27501), .ip2(\LUT[52][6] ), .op(n25927) );
  nand4_1 U29943 ( .ip1(n25930), .ip2(n25929), .ip3(n25928), .ip4(n25927), 
        .op(n25931) );
  not_ab_or_c_or_d U29944 ( .ip1(n27527), .ip2(\LUT[46][6] ), .ip3(n25932), 
        .ip4(n25931), .op(n25935) );
  nand2_1 U29945 ( .ip1(n27517), .ip2(\LUT[50][6] ), .op(n25934) );
  nand2_1 U29946 ( .ip1(n27506), .ip2(\LUT[45][6] ), .op(n25933) );
  nand4_1 U29947 ( .ip1(n25936), .ip2(n25935), .ip3(n25934), .ip4(n25933), 
        .op(n25937) );
  not_ab_or_c_or_d U29948 ( .ip1(\LUT[43][6] ), .ip2(n27519), .ip3(n25938), 
        .ip4(n25937), .op(n25939) );
  nor2_1 U29949 ( .ip1(n25939), .ip2(n27528), .op(n25945) );
  nand2_1 U29950 ( .ip1(n27563), .ip2(\LUT[62][6] ), .op(n25943) );
  nand2_1 U29951 ( .ip1(n27397), .ip2(\LUT[58][6] ), .op(n25942) );
  nand2_1 U29952 ( .ip1(n27555), .ip2(\LUT[61][6] ), .op(n25941) );
  nand2_1 U29953 ( .ip1(n27554), .ip2(\LUT[60][6] ), .op(n25940) );
  nand4_1 U29954 ( .ip1(n25943), .ip2(n25942), .ip3(n25941), .ip4(n25940), 
        .op(n25944) );
  not_ab_or_c_or_d U29955 ( .ip1(n27533), .ip2(n25946), .ip3(n25945), .ip4(
        n25944), .op(n25949) );
  nand2_1 U29956 ( .ip1(n27553), .ip2(\LUT[57][6] ), .op(n25948) );
  nand2_1 U29957 ( .ip1(n27546), .ip2(\LUT[59][6] ), .op(n25947) );
  nand4_1 U29958 ( .ip1(n25950), .ip2(n25949), .ip3(n25948), .ip4(n25947), 
        .op(n25951) );
  nand2_1 U29959 ( .ip1(n25951), .ip2(n27567), .op(n25954) );
  nand2_1 U29960 ( .ip1(n27569), .ip2(\LUT[73][6] ), .op(n25953) );
  nand2_1 U29961 ( .ip1(n27570), .ip2(\LUT[72][6] ), .op(n25952) );
  nand3_1 U29962 ( .ip1(n25954), .ip2(n25953), .ip3(n25952), .op(n25955) );
  not_ab_or_c_or_d U29963 ( .ip1(n27576), .ip2(\LUT[71][6] ), .ip3(n25956), 
        .ip4(n25955), .op(n25957) );
  inv_1 U29964 ( .ip(n27288), .op(n27577) );
  or2_1 U29965 ( .ip1(n25957), .ip2(n27577), .op(n25960) );
  nand2_1 U29966 ( .ip1(n27581), .ip2(\LUT[106][6] ), .op(n25959) );
  nand2_1 U29967 ( .ip1(n27172), .ip2(\LUT[111][6] ), .op(n25958) );
  nand4_1 U29968 ( .ip1(n25961), .ip2(n25960), .ip3(n25959), .ip4(n25958), 
        .op(n25962) );
  nand2_1 U29969 ( .ip1(n27589), .ip2(n25962), .op(n25964) );
  nand2_1 U29970 ( .ip1(sig_out[6]), .ip2(n27590), .op(n25963) );
  nand2_1 U29971 ( .ip1(n25964), .ip2(n25963), .op(n13459) );
  inv_1 U29972 ( .ip(n25965), .op(n26320) );
  and2_1 U29973 ( .ip1(n26320), .ip2(\LUT[106][7] ), .op(n25971) );
  nand2_1 U29974 ( .ip1(n27319), .ip2(\LUT[104][7] ), .op(n25969) );
  nand2_1 U29975 ( .ip1(n27318), .ip2(\LUT[107][7] ), .op(n25968) );
  nand2_1 U29976 ( .ip1(n27325), .ip2(\LUT[110][7] ), .op(n25967) );
  nand2_1 U29977 ( .ip1(n27309), .ip2(\LUT[109][7] ), .op(n25966) );
  nand4_1 U29978 ( .ip1(n25969), .ip2(n25968), .ip3(n25967), .ip4(n25966), 
        .op(n25970) );
  not_ab_or_c_or_d U29979 ( .ip1(\LUT[105][7] ), .ip2(n27317), .ip3(n25971), 
        .ip4(n25970), .op(n25975) );
  nand2_1 U29980 ( .ip1(n27328), .ip2(\LUT[101][7] ), .op(n25974) );
  nand2_1 U29981 ( .ip1(n27327), .ip2(\LUT[103][7] ), .op(n25973) );
  nand2_1 U29982 ( .ip1(n27326), .ip2(\LUT[102][7] ), .op(n25972) );
  nand4_1 U29983 ( .ip1(n25975), .ip2(n25974), .ip3(n25973), .ip4(n25972), 
        .op(n25996) );
  nand2_1 U29984 ( .ip1(n27333), .ip2(\LUT[95][7] ), .op(n25979) );
  nand2_1 U29985 ( .ip1(n27334), .ip2(\LUT[94][7] ), .op(n25978) );
  nand2_1 U29986 ( .ip1(n27335), .ip2(\LUT[98][7] ), .op(n25977) );
  nand2_1 U29987 ( .ip1(n27336), .ip2(\LUT[97][7] ), .op(n25976) );
  nand4_1 U29988 ( .ip1(n25979), .ip2(n25978), .ip3(n25977), .ip4(n25976), 
        .op(n25984) );
  nand2_1 U29989 ( .ip1(n27341), .ip2(\LUT[93][7] ), .op(n25982) );
  nand2_1 U29990 ( .ip1(n27342), .ip2(\LUT[92][7] ), .op(n25981) );
  nand2_1 U29991 ( .ip1(n27343), .ip2(\LUT[91][7] ), .op(n25980) );
  nand3_1 U29992 ( .ip1(n25982), .ip2(n25981), .ip3(n25980), .op(n25983) );
  not_ab_or_c_or_d U29993 ( .ip1(n27349), .ip2(\LUT[96][7] ), .ip3(n25984), 
        .ip4(n25983), .op(n25988) );
  nand2_1 U29994 ( .ip1(n27350), .ip2(\LUT[89][7] ), .op(n25987) );
  nand2_1 U29995 ( .ip1(n27351), .ip2(\LUT[90][7] ), .op(n25986) );
  nand2_1 U29996 ( .ip1(n27352), .ip2(\LUT[88][7] ), .op(n25985) );
  nand4_1 U29997 ( .ip1(n25988), .ip2(n25987), .ip3(n25986), .ip4(n25985), 
        .op(n25992) );
  nand2_1 U29998 ( .ip1(\LUT[85][7] ), .ip2(n27357), .op(n25990) );
  nand2_1 U29999 ( .ip1(\LUT[86][7] ), .ip2(n27358), .op(n25989) );
  nand2_1 U30000 ( .ip1(n25990), .ip2(n25989), .op(n25991) );
  not_ab_or_c_or_d U30001 ( .ip1(n27363), .ip2(\LUT[87][7] ), .ip3(n25992), 
        .ip4(n25991), .op(n25994) );
  nor2_1 U30002 ( .ip1(\LUT[99][7] ), .ip2(n27367), .op(n25993) );
  not_ab_or_c_or_d U30003 ( .ip1(n27367), .ip2(n25994), .ip3(n25993), .ip4(
        n27364), .op(n25995) );
  not_ab_or_c_or_d U30004 ( .ip1(n27370), .ip2(\LUT[100][7] ), .ip3(n25996), 
        .ip4(n25995), .op(n25997) );
  nor2_1 U30005 ( .ip1(n25997), .ip2(n27371), .op(n26007) );
  nand2_1 U30006 ( .ip1(n27298), .ip2(\LUT[117][7] ), .op(n26001) );
  nand2_1 U30007 ( .ip1(n27582), .ip2(\LUT[115][7] ), .op(n26000) );
  nand2_1 U30008 ( .ip1(n27299), .ip2(\LUT[118][7] ), .op(n25999) );
  nand2_1 U30009 ( .ip1(n27300), .ip2(\LUT[119][7] ), .op(n25998) );
  and4_1 U30010 ( .ip1(n26001), .ip2(n26000), .ip3(n25999), .ip4(n25998), .op(
        n26005) );
  nand2_1 U30011 ( .ip1(n27583), .ip2(\LUT[113][7] ), .op(n26004) );
  nand2_1 U30012 ( .ip1(n27305), .ip2(\LUT[114][7] ), .op(n26003) );
  nand2_1 U30013 ( .ip1(n27297), .ip2(\LUT[116][7] ), .op(n26002) );
  nand4_1 U30014 ( .ip1(n26005), .ip2(n26004), .ip3(n26003), .ip4(n26002), 
        .op(n26006) );
  not_ab_or_c_or_d U30015 ( .ip1(n27172), .ip2(\LUT[111][7] ), .ip3(n26007), 
        .ip4(n26006), .op(n26125) );
  and2_1 U30016 ( .ip1(n27548), .ip2(\LUT[67][7] ), .op(n26013) );
  nand2_1 U30017 ( .ip1(n27534), .ip2(\LUT[65][7] ), .op(n26011) );
  nand2_1 U30018 ( .ip1(n27537), .ip2(\LUT[68][7] ), .op(n26010) );
  nand2_1 U30019 ( .ip1(n27535), .ip2(\LUT[69][7] ), .op(n26009) );
  nand2_1 U30020 ( .ip1(n27536), .ip2(\LUT[70][7] ), .op(n26008) );
  nand4_1 U30021 ( .ip1(n26011), .ip2(n26010), .ip3(n26009), .ip4(n26008), 
        .op(n26012) );
  not_ab_or_c_or_d U30022 ( .ip1(\LUT[66][7] ), .ip2(n27542), .ip3(n26013), 
        .ip4(n26012), .op(n26017) );
  nand2_1 U30023 ( .ip1(n27546), .ip2(\LUT[59][7] ), .op(n26016) );
  nand2_1 U30024 ( .ip1(n27563), .ip2(\LUT[62][7] ), .op(n26015) );
  nand2_1 U30025 ( .ip1(n27547), .ip2(\LUT[64][7] ), .op(n26014) );
  nand4_1 U30026 ( .ip1(n26017), .ip2(n26016), .ip3(n26015), .ip4(n26014), 
        .op(n26023) );
  nand2_1 U30027 ( .ip1(n27397), .ip2(\LUT[58][7] ), .op(n26021) );
  nand2_1 U30028 ( .ip1(n27554), .ip2(\LUT[60][7] ), .op(n26020) );
  nand2_1 U30029 ( .ip1(n27555), .ip2(\LUT[61][7] ), .op(n26019) );
  nand2_1 U30030 ( .ip1(n27556), .ip2(\LUT[63][7] ), .op(n26018) );
  nand4_1 U30031 ( .ip1(n26021), .ip2(n26020), .ip3(n26019), .ip4(n26018), 
        .op(n26022) );
  not_ab_or_c_or_d U30032 ( .ip1(n27553), .ip2(\LUT[57][7] ), .ip3(n26023), 
        .ip4(n26022), .op(n26024) );
  or2_1 U30033 ( .ip1(n26024), .ip2(n27265), .op(n26102) );
  nand2_1 U30034 ( .ip1(\LUT[27][7] ), .ip2(n27398), .op(n26027) );
  nand2_1 U30035 ( .ip1(n27400), .ip2(\LUT[28][7] ), .op(n26026) );
  nand2_1 U30036 ( .ip1(n27405), .ip2(\LUT[25][7] ), .op(n26025) );
  nand3_1 U30037 ( .ip1(n26027), .ip2(n26026), .ip3(n26025), .op(n26032) );
  nand2_1 U30038 ( .ip1(\LUT[24][7] ), .ip2(n27404), .op(n26030) );
  nand2_1 U30039 ( .ip1(n27406), .ip2(\LUT[23][7] ), .op(n26029) );
  nand2_1 U30040 ( .ip1(n27399), .ip2(\LUT[26][7] ), .op(n26028) );
  nand3_1 U30041 ( .ip1(n26030), .ip2(n26029), .ip3(n26028), .op(n26031) );
  not_ab_or_c_or_d U30042 ( .ip1(n27459), .ip2(\LUT[17][7] ), .ip3(n26032), 
        .ip4(n26031), .op(n26061) );
  nand2_1 U30043 ( .ip1(\LUT[2][7] ), .ip2(n27413), .op(n26034) );
  nand2_1 U30044 ( .ip1(\LUT[3][7] ), .ip2(n27414), .op(n26033) );
  nand2_1 U30045 ( .ip1(n26034), .ip2(n26033), .op(n26050) );
  nand2_1 U30046 ( .ip1(n27428), .ip2(\LUT[6][7] ), .op(n26038) );
  nand2_1 U30047 ( .ip1(n27427), .ip2(\LUT[12][7] ), .op(n26037) );
  nand2_1 U30048 ( .ip1(n27420), .ip2(\LUT[13][7] ), .op(n26036) );
  nand2_1 U30049 ( .ip1(n27419), .ip2(\LUT[14][7] ), .op(n26035) );
  nand4_1 U30050 ( .ip1(n26038), .ip2(n26037), .ip3(n26036), .ip4(n26035), 
        .op(n26044) );
  nand2_1 U30051 ( .ip1(n27426), .ip2(\LUT[8][7] ), .op(n26042) );
  nand2_1 U30052 ( .ip1(n27435), .ip2(\LUT[11][7] ), .op(n26041) );
  nand2_1 U30053 ( .ip1(n27425), .ip2(\LUT[10][7] ), .op(n26040) );
  nand2_1 U30054 ( .ip1(n27417), .ip2(\LUT[7][7] ), .op(n26039) );
  nand4_1 U30055 ( .ip1(n26042), .ip2(n26041), .ip3(n26040), .ip4(n26039), 
        .op(n26043) );
  not_ab_or_c_or_d U30056 ( .ip1(n27418), .ip2(\LUT[9][7] ), .ip3(n26044), 
        .ip4(n26043), .op(n26048) );
  nand2_1 U30057 ( .ip1(n27436), .ip2(\LUT[0][7] ), .op(n26047) );
  nand2_1 U30058 ( .ip1(n27438), .ip2(\LUT[5][7] ), .op(n26046) );
  nand2_1 U30059 ( .ip1(n27437), .ip2(\LUT[4][7] ), .op(n26045) );
  nand4_1 U30060 ( .ip1(n26048), .ip2(n26047), .ip3(n26046), .ip4(n26045), 
        .op(n26049) );
  not_ab_or_c_or_d U30061 ( .ip1(n27445), .ip2(\LUT[1][7] ), .ip3(n26050), 
        .ip4(n26049), .op(n26051) );
  nor2_1 U30062 ( .ip1(n26051), .ip2(n27446), .op(n26057) );
  nand2_1 U30063 ( .ip1(n27448), .ip2(\LUT[18][7] ), .op(n26055) );
  nand2_1 U30064 ( .ip1(n27449), .ip2(\LUT[20][7] ), .op(n26054) );
  nand2_1 U30065 ( .ip1(n27450), .ip2(\LUT[21][7] ), .op(n26053) );
  nand2_1 U30066 ( .ip1(n27451), .ip2(\LUT[16][7] ), .op(n26052) );
  nand4_1 U30067 ( .ip1(n26055), .ip2(n26054), .ip3(n26053), .ip4(n26052), 
        .op(n26056) );
  not_ab_or_c_or_d U30068 ( .ip1(\LUT[15][7] ), .ip2(n27458), .ip3(n26057), 
        .ip4(n26056), .op(n26060) );
  nand2_1 U30069 ( .ip1(n27412), .ip2(\LUT[22][7] ), .op(n26059) );
  nand2_1 U30070 ( .ip1(n27460), .ip2(\LUT[19][7] ), .op(n26058) );
  nand4_1 U30071 ( .ip1(n26061), .ip2(n26060), .ip3(n26059), .ip4(n26058), 
        .op(n26099) );
  nand2_1 U30072 ( .ip1(\LUT[31][7] ), .ip2(n27465), .op(n26063) );
  nand2_1 U30073 ( .ip1(\LUT[30][7] ), .ip2(n27466), .op(n26062) );
  nand2_1 U30074 ( .ip1(n26063), .ip2(n26062), .op(n26078) );
  nand2_1 U30075 ( .ip1(n27470), .ip2(\LUT[38][7] ), .op(n26067) );
  nand2_1 U30076 ( .ip1(n27469), .ip2(\LUT[39][7] ), .op(n26066) );
  nand2_1 U30077 ( .ip1(n27472), .ip2(\LUT[42][7] ), .op(n26065) );
  nand2_1 U30078 ( .ip1(n27471), .ip2(\LUT[41][7] ), .op(n26064) );
  nand4_1 U30079 ( .ip1(n26067), .ip2(n26066), .ip3(n26065), .ip4(n26064), 
        .op(n26072) );
  nand2_1 U30080 ( .ip1(\LUT[36][7] ), .ip2(n27477), .op(n26070) );
  nand2_1 U30081 ( .ip1(n27478), .ip2(\LUT[37][7] ), .op(n26069) );
  nand2_1 U30082 ( .ip1(n27479), .ip2(\LUT[32][7] ), .op(n26068) );
  nand3_1 U30083 ( .ip1(n26070), .ip2(n26069), .ip3(n26068), .op(n26071) );
  not_ab_or_c_or_d U30084 ( .ip1(n27485), .ip2(\LUT[40][7] ), .ip3(n26072), 
        .ip4(n26071), .op(n26076) );
  nand2_1 U30085 ( .ip1(n27486), .ip2(\LUT[34][7] ), .op(n26075) );
  nand2_1 U30086 ( .ip1(n27488), .ip2(\LUT[33][7] ), .op(n26074) );
  nand2_1 U30087 ( .ip1(n27487), .ip2(\LUT[35][7] ), .op(n26073) );
  nand4_1 U30088 ( .ip1(n26076), .ip2(n26075), .ip3(n26074), .ip4(n26073), 
        .op(n26077) );
  not_ab_or_c_or_d U30089 ( .ip1(n27495), .ip2(\LUT[29][7] ), .ip3(n26078), 
        .ip4(n26077), .op(n26079) );
  nor2_1 U30090 ( .ip1(n26079), .ip2(n27496), .op(n26098) );
  nand2_1 U30091 ( .ip1(n27498), .ip2(\LUT[48][7] ), .op(n26083) );
  nand2_1 U30092 ( .ip1(n27499), .ip2(\LUT[49][7] ), .op(n26082) );
  nand2_1 U30093 ( .ip1(n27507), .ip2(\LUT[54][7] ), .op(n26081) );
  nand2_1 U30094 ( .ip1(n27501), .ip2(\LUT[52][7] ), .op(n26080) );
  nand4_1 U30095 ( .ip1(n26083), .ip2(n26082), .ip3(n26081), .ip4(n26080), 
        .op(n26095) );
  and2_1 U30096 ( .ip1(n27518), .ip2(\LUT[44][7] ), .op(n26089) );
  nand2_1 U30097 ( .ip1(n27508), .ip2(\LUT[55][7] ), .op(n26087) );
  nand2_1 U30098 ( .ip1(n27510), .ip2(\LUT[51][7] ), .op(n26086) );
  nand2_1 U30099 ( .ip1(n27509), .ip2(\LUT[56][7] ), .op(n26085) );
  nand2_1 U30100 ( .ip1(n27500), .ip2(\LUT[53][7] ), .op(n26084) );
  nand4_1 U30101 ( .ip1(n26087), .ip2(n26086), .ip3(n26085), .ip4(n26084), 
        .op(n26088) );
  not_ab_or_c_or_d U30102 ( .ip1(n27517), .ip2(\LUT[50][7] ), .ip3(n26089), 
        .ip4(n26088), .op(n26093) );
  nand2_1 U30103 ( .ip1(n27506), .ip2(\LUT[45][7] ), .op(n26092) );
  nand2_1 U30104 ( .ip1(n27519), .ip2(\LUT[43][7] ), .op(n26091) );
  nand2_1 U30105 ( .ip1(n27520), .ip2(\LUT[47][7] ), .op(n26090) );
  nand4_1 U30106 ( .ip1(n26093), .ip2(n26092), .ip3(n26091), .ip4(n26090), 
        .op(n26094) );
  not_ab_or_c_or_d U30107 ( .ip1(n27527), .ip2(\LUT[46][7] ), .ip3(n26095), 
        .ip4(n26094), .op(n26096) );
  nor2_1 U30108 ( .ip1(n26096), .ip2(n27528), .op(n26097) );
  not_ab_or_c_or_d U30109 ( .ip1(n27533), .ip2(n26099), .ip3(n26098), .ip4(
        n26097), .op(n26100) );
  or2_1 U30110 ( .ip1(n26100), .ip2(n27265), .op(n26101) );
  nand2_1 U30111 ( .ip1(n26102), .ip2(n26101), .op(n26116) );
  nand2_1 U30112 ( .ip1(n27391), .ip2(\LUT[75][7] ), .op(n26114) );
  nand2_1 U30113 ( .ip1(n27373), .ip2(\LUT[82][7] ), .op(n26106) );
  nand2_1 U30114 ( .ip1(n27374), .ip2(\LUT[81][7] ), .op(n26105) );
  nand2_1 U30115 ( .ip1(n27375), .ip2(\LUT[84][7] ), .op(n26104) );
  nand2_1 U30116 ( .ip1(n27376), .ip2(\LUT[83][7] ), .op(n26103) );
  nand4_1 U30117 ( .ip1(n26106), .ip2(n26105), .ip3(n26104), .ip4(n26103), 
        .op(n26111) );
  nand2_1 U30118 ( .ip1(n27381), .ip2(\LUT[78][7] ), .op(n26109) );
  nand2_1 U30119 ( .ip1(n27382), .ip2(\LUT[79][7] ), .op(n26108) );
  nand2_1 U30120 ( .ip1(n27383), .ip2(\LUT[77][7] ), .op(n26107) );
  nand3_1 U30121 ( .ip1(n26109), .ip2(n26108), .ip3(n26107), .op(n26110) );
  not_ab_or_c_or_d U30122 ( .ip1(n27389), .ip2(\LUT[80][7] ), .ip3(n26111), 
        .ip4(n26110), .op(n26113) );
  nand2_1 U30123 ( .ip1(n27392), .ip2(\LUT[74][7] ), .op(n26112) );
  nand3_1 U30124 ( .ip1(n26114), .ip2(n26113), .ip3(n26112), .op(n26115) );
  not_ab_or_c_or_d U30125 ( .ip1(n27390), .ip2(\LUT[76][7] ), .ip3(n26116), 
        .ip4(n26115), .op(n26120) );
  nand2_1 U30126 ( .ip1(n27576), .ip2(\LUT[71][7] ), .op(n26119) );
  nand2_1 U30127 ( .ip1(n27569), .ip2(\LUT[73][7] ), .op(n26118) );
  nand2_1 U30128 ( .ip1(n27570), .ip2(\LUT[72][7] ), .op(n26117) );
  nand4_1 U30129 ( .ip1(n26120), .ip2(n26119), .ip3(n26118), .ip4(n26117), 
        .op(n26121) );
  nand2_1 U30130 ( .ip1(n27288), .ip2(n26121), .op(n26124) );
  nand2_1 U30131 ( .ip1(n27165), .ip2(\LUT[108][7] ), .op(n26123) );
  nand2_1 U30132 ( .ip1(n27289), .ip2(\LUT[112][7] ), .op(n26122) );
  nand4_1 U30133 ( .ip1(n26125), .ip2(n26124), .ip3(n26123), .ip4(n26122), 
        .op(n26126) );
  nand2_1 U30134 ( .ip1(n27589), .ip2(n26126), .op(n26128) );
  nand2_1 U30135 ( .ip1(sig_out[7]), .ip2(n27590), .op(n26127) );
  nand2_1 U30136 ( .ip1(n26128), .ip2(n26127), .op(n13458) );
  nand2_1 U30137 ( .ip1(n27590), .ip2(sig_out[8]), .op(n26298) );
  nand2_1 U30138 ( .ip1(n27582), .ip2(\LUT[115][8] ), .op(n26132) );
  nand2_1 U30139 ( .ip1(n27300), .ip2(\LUT[119][8] ), .op(n26131) );
  nand2_1 U30140 ( .ip1(n27299), .ip2(\LUT[118][8] ), .op(n26130) );
  nand2_1 U30141 ( .ip1(n27298), .ip2(\LUT[117][8] ), .op(n26129) );
  and4_1 U30142 ( .ip1(n26132), .ip2(n26131), .ip3(n26130), .ip4(n26129), .op(
        n26292) );
  nand2_1 U30143 ( .ip1(n27333), .ip2(\LUT[95][8] ), .op(n26136) );
  nand2_1 U30144 ( .ip1(n27334), .ip2(\LUT[94][8] ), .op(n26135) );
  nand2_1 U30145 ( .ip1(n27335), .ip2(\LUT[98][8] ), .op(n26134) );
  nand2_1 U30146 ( .ip1(n27336), .ip2(\LUT[97][8] ), .op(n26133) );
  nand4_1 U30147 ( .ip1(n26136), .ip2(n26135), .ip3(n26134), .ip4(n26133), 
        .op(n26141) );
  nand2_1 U30148 ( .ip1(n27341), .ip2(\LUT[93][8] ), .op(n26139) );
  nand2_1 U30149 ( .ip1(n27342), .ip2(\LUT[92][8] ), .op(n26138) );
  nand2_1 U30150 ( .ip1(n27343), .ip2(\LUT[91][8] ), .op(n26137) );
  nand3_1 U30151 ( .ip1(n26139), .ip2(n26138), .ip3(n26137), .op(n26140) );
  not_ab_or_c_or_d U30152 ( .ip1(n27349), .ip2(\LUT[96][8] ), .ip3(n26141), 
        .ip4(n26140), .op(n26145) );
  nand2_1 U30153 ( .ip1(n27350), .ip2(\LUT[89][8] ), .op(n26144) );
  nand2_1 U30154 ( .ip1(n27351), .ip2(\LUT[90][8] ), .op(n26143) );
  nand2_1 U30155 ( .ip1(n27352), .ip2(\LUT[88][8] ), .op(n26142) );
  nand4_1 U30156 ( .ip1(n26145), .ip2(n26144), .ip3(n26143), .ip4(n26142), 
        .op(n26149) );
  nand2_1 U30157 ( .ip1(\LUT[85][8] ), .ip2(n27357), .op(n26147) );
  nand2_1 U30158 ( .ip1(\LUT[86][8] ), .ip2(n27358), .op(n26146) );
  nand2_1 U30159 ( .ip1(n26147), .ip2(n26146), .op(n26148) );
  not_ab_or_c_or_d U30160 ( .ip1(n27363), .ip2(\LUT[87][8] ), .ip3(n26149), 
        .ip4(n26148), .op(n26150) );
  nor2_1 U30161 ( .ip1(n26150), .ip2(n27142), .op(n26170) );
  inv_1 U30162 ( .ip(n26151), .op(n27311) );
  and2_1 U30163 ( .ip1(n27311), .ip2(\LUT[111][8] ), .op(n26154) );
  inv_1 U30164 ( .ip(n26152), .op(n27312) );
  and2_1 U30165 ( .ip1(n27312), .ip2(\LUT[112][8] ), .op(n26153) );
  not_ab_or_c_or_d U30166 ( .ip1(\LUT[110][8] ), .ip2(n27325), .ip3(n26154), 
        .ip4(n26153), .op(n26159) );
  inv_1 U30167 ( .ip(n26155), .op(n27310) );
  nand2_1 U30168 ( .ip1(n27310), .ip2(\LUT[108][8] ), .op(n26158) );
  nand2_1 U30169 ( .ip1(n27309), .ip2(\LUT[109][8] ), .op(n26157) );
  nand2_1 U30170 ( .ip1(n27318), .ip2(\LUT[107][8] ), .op(n26156) );
  nand4_1 U30171 ( .ip1(n26159), .ip2(n26158), .ip3(n26157), .ip4(n26156), 
        .op(n26164) );
  nand2_1 U30172 ( .ip1(\LUT[105][8] ), .ip2(n27317), .op(n26162) );
  nand2_1 U30173 ( .ip1(n27319), .ip2(\LUT[104][8] ), .op(n26161) );
  nand2_1 U30174 ( .ip1(n26320), .ip2(\LUT[106][8] ), .op(n26160) );
  nand3_1 U30175 ( .ip1(n26162), .ip2(n26161), .ip3(n26160), .op(n26163) );
  not_ab_or_c_or_d U30176 ( .ip1(n27328), .ip2(\LUT[101][8] ), .ip3(n26164), 
        .ip4(n26163), .op(n26168) );
  nand2_1 U30177 ( .ip1(n27156), .ip2(\LUT[99][8] ), .op(n26167) );
  nand2_1 U30178 ( .ip1(n27327), .ip2(\LUT[103][8] ), .op(n26166) );
  nand2_1 U30179 ( .ip1(n27326), .ip2(\LUT[102][8] ), .op(n26165) );
  nand4_1 U30180 ( .ip1(n26168), .ip2(n26167), .ip3(n26166), .ip4(n26165), 
        .op(n26169) );
  not_ab_or_c_or_d U30181 ( .ip1(\LUT[100][8] ), .ip2(n27370), .ip3(n26170), 
        .ip4(n26169), .op(n26171) );
  nor2_1 U30182 ( .ip1(n26171), .ip2(n27371), .op(n26288) );
  nand2_1 U30183 ( .ip1(n27373), .ip2(\LUT[82][8] ), .op(n26175) );
  nand2_1 U30184 ( .ip1(n27374), .ip2(\LUT[81][8] ), .op(n26174) );
  nand2_1 U30185 ( .ip1(n27376), .ip2(\LUT[83][8] ), .op(n26173) );
  nand2_1 U30186 ( .ip1(n27375), .ip2(\LUT[84][8] ), .op(n26172) );
  nand4_1 U30187 ( .ip1(n26175), .ip2(n26174), .ip3(n26173), .ip4(n26172), 
        .op(n26180) );
  nand2_1 U30188 ( .ip1(n27381), .ip2(\LUT[78][8] ), .op(n26178) );
  nand2_1 U30189 ( .ip1(n27382), .ip2(\LUT[79][8] ), .op(n26177) );
  nand2_1 U30190 ( .ip1(n27383), .ip2(\LUT[77][8] ), .op(n26176) );
  nand3_1 U30191 ( .ip1(n26178), .ip2(n26177), .ip3(n26176), .op(n26179) );
  not_ab_or_c_or_d U30192 ( .ip1(n27389), .ip2(\LUT[80][8] ), .ip3(n26180), 
        .ip4(n26179), .op(n26184) );
  nand2_1 U30193 ( .ip1(n27390), .ip2(\LUT[76][8] ), .op(n26183) );
  nand2_1 U30194 ( .ip1(n27391), .ip2(\LUT[75][8] ), .op(n26182) );
  nand2_1 U30195 ( .ip1(n27392), .ip2(\LUT[74][8] ), .op(n26181) );
  nand4_1 U30196 ( .ip1(n26184), .ip2(n26183), .ip3(n26182), .ip4(n26181), 
        .op(n26285) );
  nand2_1 U30197 ( .ip1(\LUT[58][8] ), .ip2(n27397), .op(n26279) );
  nand2_1 U30198 ( .ip1(n27398), .ip2(\LUT[27][8] ), .op(n26187) );
  nand2_1 U30199 ( .ip1(n27399), .ip2(\LUT[26][8] ), .op(n26186) );
  nand2_1 U30200 ( .ip1(n27400), .ip2(\LUT[28][8] ), .op(n26185) );
  nand3_1 U30201 ( .ip1(n26187), .ip2(n26186), .ip3(n26185), .op(n26192) );
  nand2_1 U30202 ( .ip1(\LUT[24][8] ), .ip2(n27404), .op(n26190) );
  nand2_1 U30203 ( .ip1(n27405), .ip2(\LUT[25][8] ), .op(n26189) );
  nand2_1 U30204 ( .ip1(n27406), .ip2(\LUT[23][8] ), .op(n26188) );
  nand3_1 U30205 ( .ip1(n26190), .ip2(n26189), .ip3(n26188), .op(n26191) );
  not_ab_or_c_or_d U30206 ( .ip1(n27459), .ip2(\LUT[17][8] ), .ip3(n26192), 
        .ip4(n26191), .op(n26221) );
  nand2_1 U30207 ( .ip1(\LUT[2][8] ), .ip2(n27413), .op(n26194) );
  nand2_1 U30208 ( .ip1(\LUT[3][8] ), .ip2(n27414), .op(n26193) );
  nand2_1 U30209 ( .ip1(n26194), .ip2(n26193), .op(n26210) );
  nand2_1 U30210 ( .ip1(n27427), .ip2(\LUT[12][8] ), .op(n26198) );
  nand2_1 U30211 ( .ip1(n27428), .ip2(\LUT[6][8] ), .op(n26197) );
  nand2_1 U30212 ( .ip1(n27419), .ip2(\LUT[14][8] ), .op(n26196) );
  nand2_1 U30213 ( .ip1(n27420), .ip2(\LUT[13][8] ), .op(n26195) );
  nand4_1 U30214 ( .ip1(n26198), .ip2(n26197), .ip3(n26196), .ip4(n26195), 
        .op(n26204) );
  nand2_1 U30215 ( .ip1(n27425), .ip2(\LUT[10][8] ), .op(n26202) );
  nand2_1 U30216 ( .ip1(n27435), .ip2(\LUT[11][8] ), .op(n26201) );
  nand2_1 U30217 ( .ip1(n27417), .ip2(\LUT[7][8] ), .op(n26200) );
  nand2_1 U30218 ( .ip1(n27426), .ip2(\LUT[8][8] ), .op(n26199) );
  nand4_1 U30219 ( .ip1(n26202), .ip2(n26201), .ip3(n26200), .ip4(n26199), 
        .op(n26203) );
  not_ab_or_c_or_d U30220 ( .ip1(n27418), .ip2(\LUT[9][8] ), .ip3(n26204), 
        .ip4(n26203), .op(n26208) );
  nand2_1 U30221 ( .ip1(n27445), .ip2(\LUT[1][8] ), .op(n26207) );
  nand2_1 U30222 ( .ip1(n27437), .ip2(\LUT[4][8] ), .op(n26206) );
  nand2_1 U30223 ( .ip1(n27438), .ip2(\LUT[5][8] ), .op(n26205) );
  nand4_1 U30224 ( .ip1(n26208), .ip2(n26207), .ip3(n26206), .ip4(n26205), 
        .op(n26209) );
  not_ab_or_c_or_d U30225 ( .ip1(n27436), .ip2(\LUT[0][8] ), .ip3(n26210), 
        .ip4(n26209), .op(n26211) );
  nor2_1 U30226 ( .ip1(n26211), .ip2(n27446), .op(n26217) );
  nand2_1 U30227 ( .ip1(n27450), .ip2(\LUT[21][8] ), .op(n26215) );
  nand2_1 U30228 ( .ip1(n27449), .ip2(\LUT[20][8] ), .op(n26214) );
  nand2_1 U30229 ( .ip1(n27451), .ip2(\LUT[16][8] ), .op(n26213) );
  nand2_1 U30230 ( .ip1(n27448), .ip2(\LUT[18][8] ), .op(n26212) );
  nand4_1 U30231 ( .ip1(n26215), .ip2(n26214), .ip3(n26213), .ip4(n26212), 
        .op(n26216) );
  not_ab_or_c_or_d U30232 ( .ip1(\LUT[15][8] ), .ip2(n27458), .ip3(n26217), 
        .ip4(n26216), .op(n26220) );
  nand2_1 U30233 ( .ip1(n27412), .ip2(\LUT[22][8] ), .op(n26219) );
  nand2_1 U30234 ( .ip1(n27460), .ip2(\LUT[19][8] ), .op(n26218) );
  nand4_1 U30235 ( .ip1(n26221), .ip2(n26220), .ip3(n26219), .ip4(n26218), 
        .op(n26259) );
  nand2_1 U30236 ( .ip1(n27527), .ip2(\LUT[46][8] ), .op(n26225) );
  nand2_1 U30237 ( .ip1(n27498), .ip2(\LUT[48][8] ), .op(n26224) );
  nand2_1 U30238 ( .ip1(n27501), .ip2(\LUT[52][8] ), .op(n26223) );
  nand2_1 U30239 ( .ip1(n27500), .ip2(\LUT[53][8] ), .op(n26222) );
  nand4_1 U30240 ( .ip1(n26225), .ip2(n26224), .ip3(n26223), .ip4(n26222), 
        .op(n26237) );
  and2_1 U30241 ( .ip1(n27499), .ip2(\LUT[49][8] ), .op(n26231) );
  nand2_1 U30242 ( .ip1(n27507), .ip2(\LUT[54][8] ), .op(n26229) );
  nand2_1 U30243 ( .ip1(n27510), .ip2(\LUT[51][8] ), .op(n26228) );
  nand2_1 U30244 ( .ip1(n27509), .ip2(\LUT[56][8] ), .op(n26227) );
  nand2_1 U30245 ( .ip1(n27508), .ip2(\LUT[55][8] ), .op(n26226) );
  nand4_1 U30246 ( .ip1(n26229), .ip2(n26228), .ip3(n26227), .ip4(n26226), 
        .op(n26230) );
  not_ab_or_c_or_d U30247 ( .ip1(n27506), .ip2(\LUT[45][8] ), .ip3(n26231), 
        .ip4(n26230), .op(n26235) );
  nand2_1 U30248 ( .ip1(n27519), .ip2(\LUT[43][8] ), .op(n26234) );
  nand2_1 U30249 ( .ip1(n27518), .ip2(\LUT[44][8] ), .op(n26233) );
  nand2_1 U30250 ( .ip1(n27520), .ip2(\LUT[47][8] ), .op(n26232) );
  nand4_1 U30251 ( .ip1(n26235), .ip2(n26234), .ip3(n26233), .ip4(n26232), 
        .op(n26236) );
  not_ab_or_c_or_d U30252 ( .ip1(n27517), .ip2(\LUT[50][8] ), .ip3(n26237), 
        .ip4(n26236), .op(n26238) );
  nor2_1 U30253 ( .ip1(n26238), .ip2(n27528), .op(n26258) );
  nand2_1 U30254 ( .ip1(\LUT[31][8] ), .ip2(n27465), .op(n26240) );
  nand2_1 U30255 ( .ip1(\LUT[30][8] ), .ip2(n27466), .op(n26239) );
  nand2_1 U30256 ( .ip1(n26240), .ip2(n26239), .op(n26255) );
  nand2_1 U30257 ( .ip1(n27469), .ip2(\LUT[39][8] ), .op(n26244) );
  nand2_1 U30258 ( .ip1(n27470), .ip2(\LUT[38][8] ), .op(n26243) );
  nand2_1 U30259 ( .ip1(n27471), .ip2(\LUT[41][8] ), .op(n26242) );
  nand2_1 U30260 ( .ip1(n27472), .ip2(\LUT[42][8] ), .op(n26241) );
  nand4_1 U30261 ( .ip1(n26244), .ip2(n26243), .ip3(n26242), .ip4(n26241), 
        .op(n26249) );
  nand2_1 U30262 ( .ip1(\LUT[36][8] ), .ip2(n27477), .op(n26247) );
  nand2_1 U30263 ( .ip1(n27478), .ip2(\LUT[37][8] ), .op(n26246) );
  nand2_1 U30264 ( .ip1(n27479), .ip2(\LUT[32][8] ), .op(n26245) );
  nand3_1 U30265 ( .ip1(n26247), .ip2(n26246), .ip3(n26245), .op(n26248) );
  not_ab_or_c_or_d U30266 ( .ip1(n27485), .ip2(\LUT[40][8] ), .ip3(n26249), 
        .ip4(n26248), .op(n26253) );
  nand2_1 U30267 ( .ip1(n27486), .ip2(\LUT[34][8] ), .op(n26252) );
  nand2_1 U30268 ( .ip1(n27487), .ip2(\LUT[35][8] ), .op(n26251) );
  nand2_1 U30269 ( .ip1(n27488), .ip2(\LUT[33][8] ), .op(n26250) );
  nand4_1 U30270 ( .ip1(n26253), .ip2(n26252), .ip3(n26251), .ip4(n26250), 
        .op(n26254) );
  not_ab_or_c_or_d U30271 ( .ip1(n27495), .ip2(\LUT[29][8] ), .ip3(n26255), 
        .ip4(n26254), .op(n26256) );
  nor2_1 U30272 ( .ip1(n26256), .ip2(n27496), .op(n26257) );
  not_ab_or_c_or_d U30273 ( .ip1(n27533), .ip2(n26259), .ip3(n26258), .ip4(
        n26257), .op(n26278) );
  nand2_1 U30274 ( .ip1(n27534), .ip2(\LUT[65][8] ), .op(n26263) );
  nand2_1 U30275 ( .ip1(n27537), .ip2(\LUT[68][8] ), .op(n26262) );
  nand2_1 U30276 ( .ip1(n27535), .ip2(\LUT[69][8] ), .op(n26261) );
  nand2_1 U30277 ( .ip1(n27536), .ip2(\LUT[70][8] ), .op(n26260) );
  nand4_1 U30278 ( .ip1(n26263), .ip2(n26262), .ip3(n26261), .ip4(n26260), 
        .op(n26264) );
  or2_1 U30279 ( .ip1(n27548), .ip2(n26264), .op(n26266) );
  or2_1 U30280 ( .ip1(\LUT[67][8] ), .ip2(n26264), .op(n26265) );
  nand2_1 U30281 ( .ip1(n26266), .ip2(n26265), .op(n26270) );
  nand2_1 U30282 ( .ip1(n27547), .ip2(\LUT[64][8] ), .op(n26269) );
  nand2_1 U30283 ( .ip1(n27556), .ip2(\LUT[63][8] ), .op(n26268) );
  nand2_1 U30284 ( .ip1(n27542), .ip2(\LUT[66][8] ), .op(n26267) );
  nand4_1 U30285 ( .ip1(n26270), .ip2(n26269), .ip3(n26268), .ip4(n26267), 
        .op(n26276) );
  nand2_1 U30286 ( .ip1(n27553), .ip2(\LUT[57][8] ), .op(n26274) );
  nand2_1 U30287 ( .ip1(n27554), .ip2(\LUT[60][8] ), .op(n26273) );
  nand2_1 U30288 ( .ip1(n27563), .ip2(\LUT[62][8] ), .op(n26272) );
  nand2_1 U30289 ( .ip1(n27555), .ip2(\LUT[61][8] ), .op(n26271) );
  nand4_1 U30290 ( .ip1(n26274), .ip2(n26273), .ip3(n26272), .ip4(n26271), 
        .op(n26275) );
  not_ab_or_c_or_d U30291 ( .ip1(n27546), .ip2(\LUT[59][8] ), .ip3(n26276), 
        .ip4(n26275), .op(n26277) );
  nand3_1 U30292 ( .ip1(n26279), .ip2(n26278), .ip3(n26277), .op(n26280) );
  nand2_1 U30293 ( .ip1(n26280), .ip2(n27567), .op(n26283) );
  nand2_1 U30294 ( .ip1(n27569), .ip2(\LUT[73][8] ), .op(n26282) );
  nand2_1 U30295 ( .ip1(n27570), .ip2(\LUT[72][8] ), .op(n26281) );
  nand3_1 U30296 ( .ip1(n26283), .ip2(n26282), .ip3(n26281), .op(n26284) );
  not_ab_or_c_or_d U30297 ( .ip1(n27576), .ip2(\LUT[71][8] ), .ip3(n26285), 
        .ip4(n26284), .op(n26286) );
  nor2_1 U30298 ( .ip1(n26286), .ip2(n27577), .op(n26287) );
  not_ab_or_c_or_d U30299 ( .ip1(n27583), .ip2(\LUT[113][8] ), .ip3(n26288), 
        .ip4(n26287), .op(n26291) );
  nand2_1 U30300 ( .ip1(n27297), .ip2(\LUT[116][8] ), .op(n26290) );
  nand2_1 U30301 ( .ip1(n27305), .ip2(\LUT[114][8] ), .op(n26289) );
  nand4_1 U30302 ( .ip1(n26292), .ip2(n26291), .ip3(n26290), .ip4(n26289), 
        .op(n26293) );
  nand2_1 U30303 ( .ip1(n27589), .ip2(n26293), .op(n26297) );
  nand2_1 U30304 ( .ip1(n26295), .ip2(n26294), .op(n26296) );
  nand3_1 U30305 ( .ip1(n26298), .ip2(n26297), .ip3(n26296), .op(n13457) );
  nand2_1 U30306 ( .ip1(n27333), .ip2(\LUT[95][9] ), .op(n26302) );
  nand2_1 U30307 ( .ip1(n27334), .ip2(\LUT[94][9] ), .op(n26301) );
  nand2_1 U30308 ( .ip1(n27335), .ip2(\LUT[98][9] ), .op(n26300) );
  nand2_1 U30309 ( .ip1(n27336), .ip2(\LUT[97][9] ), .op(n26299) );
  nand4_1 U30310 ( .ip1(n26302), .ip2(n26301), .ip3(n26300), .ip4(n26299), 
        .op(n26307) );
  nand2_1 U30311 ( .ip1(n27341), .ip2(\LUT[93][9] ), .op(n26305) );
  nand2_1 U30312 ( .ip1(n27342), .ip2(\LUT[92][9] ), .op(n26304) );
  nand2_1 U30313 ( .ip1(n27343), .ip2(\LUT[91][9] ), .op(n26303) );
  nand3_1 U30314 ( .ip1(n26305), .ip2(n26304), .ip3(n26303), .op(n26306) );
  not_ab_or_c_or_d U30315 ( .ip1(n27349), .ip2(\LUT[96][9] ), .ip3(n26307), 
        .ip4(n26306), .op(n26311) );
  nand2_1 U30316 ( .ip1(n27350), .ip2(\LUT[89][9] ), .op(n26310) );
  nand2_1 U30317 ( .ip1(n27351), .ip2(\LUT[90][9] ), .op(n26309) );
  nand2_1 U30318 ( .ip1(n27352), .ip2(\LUT[88][9] ), .op(n26308) );
  nand4_1 U30319 ( .ip1(n26311), .ip2(n26310), .ip3(n26309), .ip4(n26308), 
        .op(n26315) );
  nand2_1 U30320 ( .ip1(\LUT[85][9] ), .ip2(n27357), .op(n26313) );
  nand2_1 U30321 ( .ip1(\LUT[86][9] ), .ip2(n27358), .op(n26312) );
  nand2_1 U30322 ( .ip1(n26313), .ip2(n26312), .op(n26314) );
  not_ab_or_c_or_d U30323 ( .ip1(n27363), .ip2(\LUT[87][9] ), .ip3(n26315), 
        .ip4(n26314), .op(n26316) );
  nor2_1 U30324 ( .ip1(n26316), .ip2(n27142), .op(n26331) );
  nand2_1 U30325 ( .ip1(n27318), .ip2(\LUT[107][9] ), .op(n26319) );
  nand2_1 U30326 ( .ip1(n27309), .ip2(\LUT[109][9] ), .op(n26318) );
  nand2_1 U30327 ( .ip1(n27325), .ip2(\LUT[110][9] ), .op(n26317) );
  nand3_1 U30328 ( .ip1(n26319), .ip2(n26318), .ip3(n26317), .op(n26325) );
  nand2_1 U30329 ( .ip1(n27317), .ip2(\LUT[105][9] ), .op(n26323) );
  nand2_1 U30330 ( .ip1(n26320), .ip2(\LUT[106][9] ), .op(n26322) );
  nand2_1 U30331 ( .ip1(n27319), .ip2(\LUT[104][9] ), .op(n26321) );
  nand3_1 U30332 ( .ip1(n26323), .ip2(n26322), .ip3(n26321), .op(n26324) );
  not_ab_or_c_or_d U30333 ( .ip1(n27326), .ip2(\LUT[102][9] ), .ip3(n26325), 
        .ip4(n26324), .op(n26329) );
  nand2_1 U30334 ( .ip1(n27370), .ip2(\LUT[100][9] ), .op(n26328) );
  nand2_1 U30335 ( .ip1(n27328), .ip2(\LUT[101][9] ), .op(n26327) );
  nand2_1 U30336 ( .ip1(n27327), .ip2(\LUT[103][9] ), .op(n26326) );
  nand4_1 U30337 ( .ip1(n26329), .ip2(n26328), .ip3(n26327), .ip4(n26326), 
        .op(n26330) );
  not_ab_or_c_or_d U30338 ( .ip1(\LUT[99][9] ), .ip2(n27156), .ip3(n26331), 
        .ip4(n26330), .op(n26332) );
  nor2_1 U30339 ( .ip1(n26332), .ip2(n27371), .op(n26342) );
  nand2_1 U30340 ( .ip1(n27298), .ip2(\LUT[117][9] ), .op(n26336) );
  nand2_1 U30341 ( .ip1(n27582), .ip2(\LUT[115][9] ), .op(n26335) );
  nand2_1 U30342 ( .ip1(n27299), .ip2(\LUT[118][9] ), .op(n26334) );
  nand2_1 U30343 ( .ip1(n27300), .ip2(\LUT[119][9] ), .op(n26333) );
  and4_1 U30344 ( .ip1(n26336), .ip2(n26335), .ip3(n26334), .ip4(n26333), .op(
        n26340) );
  nand2_1 U30345 ( .ip1(n27583), .ip2(\LUT[113][9] ), .op(n26339) );
  nand2_1 U30346 ( .ip1(n27305), .ip2(\LUT[114][9] ), .op(n26338) );
  nand2_1 U30347 ( .ip1(n27297), .ip2(\LUT[116][9] ), .op(n26337) );
  nand4_1 U30348 ( .ip1(n26340), .ip2(n26339), .ip3(n26338), .ip4(n26337), 
        .op(n26341) );
  not_ab_or_c_or_d U30349 ( .ip1(n27172), .ip2(\LUT[111][9] ), .ip3(n26342), 
        .ip4(n26341), .op(n26460) );
  and2_1 U30350 ( .ip1(n27534), .ip2(\LUT[65][9] ), .op(n26348) );
  nand2_1 U30351 ( .ip1(n27548), .ip2(\LUT[67][9] ), .op(n26346) );
  nand2_1 U30352 ( .ip1(n27537), .ip2(\LUT[68][9] ), .op(n26345) );
  nand2_1 U30353 ( .ip1(n27536), .ip2(\LUT[70][9] ), .op(n26344) );
  nand2_1 U30354 ( .ip1(n27535), .ip2(\LUT[69][9] ), .op(n26343) );
  nand4_1 U30355 ( .ip1(n26346), .ip2(n26345), .ip3(n26344), .ip4(n26343), 
        .op(n26347) );
  not_ab_or_c_or_d U30356 ( .ip1(n27542), .ip2(\LUT[66][9] ), .ip3(n26348), 
        .ip4(n26347), .op(n26352) );
  nand2_1 U30357 ( .ip1(n27547), .ip2(\LUT[64][9] ), .op(n26351) );
  nand2_1 U30358 ( .ip1(n27546), .ip2(\LUT[59][9] ), .op(n26350) );
  nand2_1 U30359 ( .ip1(n27555), .ip2(\LUT[61][9] ), .op(n26349) );
  nand4_1 U30360 ( .ip1(n26352), .ip2(n26351), .ip3(n26350), .ip4(n26349), 
        .op(n26358) );
  nand2_1 U30361 ( .ip1(n27397), .ip2(\LUT[58][9] ), .op(n26356) );
  nand2_1 U30362 ( .ip1(n27563), .ip2(\LUT[62][9] ), .op(n26355) );
  nand2_1 U30363 ( .ip1(n27556), .ip2(\LUT[63][9] ), .op(n26354) );
  nand2_1 U30364 ( .ip1(n27554), .ip2(\LUT[60][9] ), .op(n26353) );
  nand4_1 U30365 ( .ip1(n26356), .ip2(n26355), .ip3(n26354), .ip4(n26353), 
        .op(n26357) );
  not_ab_or_c_or_d U30366 ( .ip1(n27553), .ip2(\LUT[57][9] ), .ip3(n26358), 
        .ip4(n26357), .op(n26359) );
  or2_1 U30367 ( .ip1(n26359), .ip2(n27265), .op(n26437) );
  nand2_1 U30368 ( .ip1(\LUT[27][9] ), .ip2(n27398), .op(n26362) );
  nand2_1 U30369 ( .ip1(n27405), .ip2(\LUT[25][9] ), .op(n26361) );
  nand2_1 U30370 ( .ip1(n27400), .ip2(\LUT[28][9] ), .op(n26360) );
  nand3_1 U30371 ( .ip1(n26362), .ip2(n26361), .ip3(n26360), .op(n26367) );
  nand2_1 U30372 ( .ip1(\LUT[24][9] ), .ip2(n27404), .op(n26365) );
  nand2_1 U30373 ( .ip1(n27399), .ip2(\LUT[26][9] ), .op(n26364) );
  nand2_1 U30374 ( .ip1(n27406), .ip2(\LUT[23][9] ), .op(n26363) );
  nand3_1 U30375 ( .ip1(n26365), .ip2(n26364), .ip3(n26363), .op(n26366) );
  not_ab_or_c_or_d U30376 ( .ip1(n27460), .ip2(\LUT[19][9] ), .ip3(n26367), 
        .ip4(n26366), .op(n26396) );
  nand2_1 U30377 ( .ip1(\LUT[2][9] ), .ip2(n27413), .op(n26369) );
  nand2_1 U30378 ( .ip1(\LUT[3][9] ), .ip2(n27414), .op(n26368) );
  nand2_1 U30379 ( .ip1(n26369), .ip2(n26368), .op(n26385) );
  nand2_1 U30380 ( .ip1(n27427), .ip2(\LUT[12][9] ), .op(n26373) );
  nand2_1 U30381 ( .ip1(n27428), .ip2(\LUT[6][9] ), .op(n26372) );
  nand2_1 U30382 ( .ip1(n27419), .ip2(\LUT[14][9] ), .op(n26371) );
  nand2_1 U30383 ( .ip1(n27420), .ip2(\LUT[13][9] ), .op(n26370) );
  nand4_1 U30384 ( .ip1(n26373), .ip2(n26372), .ip3(n26371), .ip4(n26370), 
        .op(n26379) );
  nand2_1 U30385 ( .ip1(n27435), .ip2(\LUT[11][9] ), .op(n26377) );
  nand2_1 U30386 ( .ip1(n27425), .ip2(\LUT[10][9] ), .op(n26376) );
  nand2_1 U30387 ( .ip1(n27426), .ip2(\LUT[8][9] ), .op(n26375) );
  nand2_1 U30388 ( .ip1(n27417), .ip2(\LUT[7][9] ), .op(n26374) );
  nand4_1 U30389 ( .ip1(n26377), .ip2(n26376), .ip3(n26375), .ip4(n26374), 
        .op(n26378) );
  not_ab_or_c_or_d U30390 ( .ip1(n27418), .ip2(\LUT[9][9] ), .ip3(n26379), 
        .ip4(n26378), .op(n26383) );
  nand2_1 U30391 ( .ip1(n27436), .ip2(\LUT[0][9] ), .op(n26382) );
  nand2_1 U30392 ( .ip1(n27438), .ip2(\LUT[5][9] ), .op(n26381) );
  nand2_1 U30393 ( .ip1(n27437), .ip2(\LUT[4][9] ), .op(n26380) );
  nand4_1 U30394 ( .ip1(n26383), .ip2(n26382), .ip3(n26381), .ip4(n26380), 
        .op(n26384) );
  not_ab_or_c_or_d U30395 ( .ip1(n27445), .ip2(\LUT[1][9] ), .ip3(n26385), 
        .ip4(n26384), .op(n26386) );
  nor2_1 U30396 ( .ip1(n26386), .ip2(n27446), .op(n26392) );
  nand2_1 U30397 ( .ip1(n27450), .ip2(\LUT[21][9] ), .op(n26390) );
  nand2_1 U30398 ( .ip1(n27451), .ip2(\LUT[16][9] ), .op(n26389) );
  nand2_1 U30399 ( .ip1(n27448), .ip2(\LUT[18][9] ), .op(n26388) );
  nand2_1 U30400 ( .ip1(n27449), .ip2(\LUT[20][9] ), .op(n26387) );
  nand4_1 U30401 ( .ip1(n26390), .ip2(n26389), .ip3(n26388), .ip4(n26387), 
        .op(n26391) );
  not_ab_or_c_or_d U30402 ( .ip1(\LUT[15][9] ), .ip2(n27458), .ip3(n26392), 
        .ip4(n26391), .op(n26395) );
  nand2_1 U30403 ( .ip1(n27412), .ip2(\LUT[22][9] ), .op(n26394) );
  nand2_1 U30404 ( .ip1(n27459), .ip2(\LUT[17][9] ), .op(n26393) );
  nand4_1 U30405 ( .ip1(n26396), .ip2(n26395), .ip3(n26394), .ip4(n26393), 
        .op(n26434) );
  nand2_1 U30406 ( .ip1(\LUT[31][9] ), .ip2(n27465), .op(n26398) );
  nand2_1 U30407 ( .ip1(\LUT[30][9] ), .ip2(n27466), .op(n26397) );
  nand2_1 U30408 ( .ip1(n26398), .ip2(n26397), .op(n26413) );
  nand2_1 U30409 ( .ip1(n27469), .ip2(\LUT[39][9] ), .op(n26402) );
  nand2_1 U30410 ( .ip1(n27470), .ip2(\LUT[38][9] ), .op(n26401) );
  nand2_1 U30411 ( .ip1(n27471), .ip2(\LUT[41][9] ), .op(n26400) );
  nand2_1 U30412 ( .ip1(n27472), .ip2(\LUT[42][9] ), .op(n26399) );
  nand4_1 U30413 ( .ip1(n26402), .ip2(n26401), .ip3(n26400), .ip4(n26399), 
        .op(n26407) );
  nand2_1 U30414 ( .ip1(\LUT[36][9] ), .ip2(n27477), .op(n26405) );
  nand2_1 U30415 ( .ip1(n27478), .ip2(\LUT[37][9] ), .op(n26404) );
  nand2_1 U30416 ( .ip1(n27488), .ip2(\LUT[33][9] ), .op(n26403) );
  nand3_1 U30417 ( .ip1(n26405), .ip2(n26404), .ip3(n26403), .op(n26406) );
  not_ab_or_c_or_d U30418 ( .ip1(n27485), .ip2(\LUT[40][9] ), .ip3(n26407), 
        .ip4(n26406), .op(n26411) );
  nand2_1 U30419 ( .ip1(n27487), .ip2(\LUT[35][9] ), .op(n26410) );
  nand2_1 U30420 ( .ip1(n27486), .ip2(\LUT[34][9] ), .op(n26409) );
  nand2_1 U30421 ( .ip1(n27479), .ip2(\LUT[32][9] ), .op(n26408) );
  nand4_1 U30422 ( .ip1(n26411), .ip2(n26410), .ip3(n26409), .ip4(n26408), 
        .op(n26412) );
  not_ab_or_c_or_d U30423 ( .ip1(n27495), .ip2(\LUT[29][9] ), .ip3(n26413), 
        .ip4(n26412), .op(n26414) );
  nor2_1 U30424 ( .ip1(n26414), .ip2(n27496), .op(n26433) );
  nand2_1 U30425 ( .ip1(n27527), .ip2(\LUT[46][9] ), .op(n26418) );
  nand2_1 U30426 ( .ip1(n27498), .ip2(\LUT[48][9] ), .op(n26417) );
  nand2_1 U30427 ( .ip1(n27501), .ip2(\LUT[52][9] ), .op(n26416) );
  nand2_1 U30428 ( .ip1(n27500), .ip2(\LUT[53][9] ), .op(n26415) );
  nand4_1 U30429 ( .ip1(n26418), .ip2(n26417), .ip3(n26416), .ip4(n26415), 
        .op(n26430) );
  and2_1 U30430 ( .ip1(n27499), .ip2(\LUT[49][9] ), .op(n26424) );
  nand2_1 U30431 ( .ip1(n27507), .ip2(\LUT[54][9] ), .op(n26422) );
  nand2_1 U30432 ( .ip1(n27510), .ip2(\LUT[51][9] ), .op(n26421) );
  nand2_1 U30433 ( .ip1(n27509), .ip2(\LUT[56][9] ), .op(n26420) );
  nand2_1 U30434 ( .ip1(n27508), .ip2(\LUT[55][9] ), .op(n26419) );
  nand4_1 U30435 ( .ip1(n26422), .ip2(n26421), .ip3(n26420), .ip4(n26419), 
        .op(n26423) );
  not_ab_or_c_or_d U30436 ( .ip1(\LUT[45][9] ), .ip2(n27506), .ip3(n26424), 
        .ip4(n26423), .op(n26428) );
  nand2_1 U30437 ( .ip1(n27519), .ip2(\LUT[43][9] ), .op(n26427) );
  nand2_1 U30438 ( .ip1(n27518), .ip2(\LUT[44][9] ), .op(n26426) );
  nand2_1 U30439 ( .ip1(n27520), .ip2(\LUT[47][9] ), .op(n26425) );
  nand4_1 U30440 ( .ip1(n26428), .ip2(n26427), .ip3(n26426), .ip4(n26425), 
        .op(n26429) );
  not_ab_or_c_or_d U30441 ( .ip1(n27517), .ip2(\LUT[50][9] ), .ip3(n26430), 
        .ip4(n26429), .op(n26431) );
  nor2_1 U30442 ( .ip1(n26431), .ip2(n27528), .op(n26432) );
  not_ab_or_c_or_d U30443 ( .ip1(n27533), .ip2(n26434), .ip3(n26433), .ip4(
        n26432), .op(n26435) );
  or2_1 U30444 ( .ip1(n26435), .ip2(n27265), .op(n26436) );
  nand2_1 U30445 ( .ip1(n26437), .ip2(n26436), .op(n26451) );
  nand2_1 U30446 ( .ip1(n27391), .ip2(\LUT[75][9] ), .op(n26449) );
  nand2_1 U30447 ( .ip1(n27373), .ip2(\LUT[82][9] ), .op(n26441) );
  nand2_1 U30448 ( .ip1(n27374), .ip2(\LUT[81][9] ), .op(n26440) );
  nand2_1 U30449 ( .ip1(n27376), .ip2(\LUT[83][9] ), .op(n26439) );
  nand2_1 U30450 ( .ip1(n27375), .ip2(\LUT[84][9] ), .op(n26438) );
  nand4_1 U30451 ( .ip1(n26441), .ip2(n26440), .ip3(n26439), .ip4(n26438), 
        .op(n26446) );
  nand2_1 U30452 ( .ip1(n27381), .ip2(\LUT[78][9] ), .op(n26444) );
  nand2_1 U30453 ( .ip1(n27382), .ip2(\LUT[79][9] ), .op(n26443) );
  nand2_1 U30454 ( .ip1(n27383), .ip2(\LUT[77][9] ), .op(n26442) );
  nand3_1 U30455 ( .ip1(n26444), .ip2(n26443), .ip3(n26442), .op(n26445) );
  not_ab_or_c_or_d U30456 ( .ip1(n27389), .ip2(\LUT[80][9] ), .ip3(n26446), 
        .ip4(n26445), .op(n26448) );
  nand2_1 U30457 ( .ip1(n27392), .ip2(\LUT[74][9] ), .op(n26447) );
  nand3_1 U30458 ( .ip1(n26449), .ip2(n26448), .ip3(n26447), .op(n26450) );
  not_ab_or_c_or_d U30459 ( .ip1(n27390), .ip2(\LUT[76][9] ), .ip3(n26451), 
        .ip4(n26450), .op(n26455) );
  nand2_1 U30460 ( .ip1(n27576), .ip2(\LUT[71][9] ), .op(n26454) );
  nand2_1 U30461 ( .ip1(n27569), .ip2(\LUT[73][9] ), .op(n26453) );
  nand2_1 U30462 ( .ip1(n27570), .ip2(\LUT[72][9] ), .op(n26452) );
  nand4_1 U30463 ( .ip1(n26455), .ip2(n26454), .ip3(n26453), .ip4(n26452), 
        .op(n26456) );
  nand2_1 U30464 ( .ip1(n27288), .ip2(n26456), .op(n26459) );
  nand2_1 U30465 ( .ip1(n27165), .ip2(\LUT[108][9] ), .op(n26458) );
  nand2_1 U30466 ( .ip1(n27289), .ip2(\LUT[112][9] ), .op(n26457) );
  nand4_1 U30467 ( .ip1(n26460), .ip2(n26459), .ip3(n26458), .ip4(n26457), 
        .op(n26461) );
  nand2_1 U30468 ( .ip1(n27589), .ip2(n26461), .op(n26463) );
  nand2_1 U30469 ( .ip1(sig_out[9]), .ip2(n27590), .op(n26462) );
  nand2_1 U30470 ( .ip1(n26463), .ip2(n26462), .op(n13456) );
  nand2_1 U30471 ( .ip1(n27333), .ip2(\LUT[95][10] ), .op(n26467) );
  nand2_1 U30472 ( .ip1(n27334), .ip2(\LUT[94][10] ), .op(n26466) );
  nand2_1 U30473 ( .ip1(n27336), .ip2(\LUT[97][10] ), .op(n26465) );
  nand2_1 U30474 ( .ip1(n27335), .ip2(\LUT[98][10] ), .op(n26464) );
  nand4_1 U30475 ( .ip1(n26467), .ip2(n26466), .ip3(n26465), .ip4(n26464), 
        .op(n26472) );
  nand2_1 U30476 ( .ip1(n27341), .ip2(\LUT[93][10] ), .op(n26470) );
  nand2_1 U30477 ( .ip1(n27342), .ip2(\LUT[92][10] ), .op(n26469) );
  nand2_1 U30478 ( .ip1(n27343), .ip2(\LUT[91][10] ), .op(n26468) );
  nand3_1 U30479 ( .ip1(n26470), .ip2(n26469), .ip3(n26468), .op(n26471) );
  not_ab_or_c_or_d U30480 ( .ip1(n27349), .ip2(\LUT[96][10] ), .ip3(n26472), 
        .ip4(n26471), .op(n26476) );
  nand2_1 U30481 ( .ip1(n27350), .ip2(\LUT[89][10] ), .op(n26475) );
  nand2_1 U30482 ( .ip1(n27351), .ip2(\LUT[90][10] ), .op(n26474) );
  nand2_1 U30483 ( .ip1(n27352), .ip2(\LUT[88][10] ), .op(n26473) );
  nand4_1 U30484 ( .ip1(n26476), .ip2(n26475), .ip3(n26474), .ip4(n26473), 
        .op(n26480) );
  nand2_1 U30485 ( .ip1(\LUT[85][10] ), .ip2(n27357), .op(n26478) );
  nand2_1 U30486 ( .ip1(\LUT[86][10] ), .ip2(n27358), .op(n26477) );
  nand2_1 U30487 ( .ip1(n26478), .ip2(n26477), .op(n26479) );
  not_ab_or_c_or_d U30488 ( .ip1(n27363), .ip2(\LUT[87][10] ), .ip3(n26480), 
        .ip4(n26479), .op(n26481) );
  nor2_1 U30489 ( .ip1(n26481), .ip2(n27142), .op(n26493) );
  and2_1 U30490 ( .ip1(n27317), .ip2(\LUT[105][10] ), .op(n26487) );
  nand2_1 U30491 ( .ip1(n27318), .ip2(\LUT[107][10] ), .op(n26485) );
  nand2_1 U30492 ( .ip1(n27319), .ip2(\LUT[104][10] ), .op(n26484) );
  nand2_1 U30493 ( .ip1(n27309), .ip2(\LUT[109][10] ), .op(n26483) );
  nand2_1 U30494 ( .ip1(n27325), .ip2(\LUT[110][10] ), .op(n26482) );
  nand4_1 U30495 ( .ip1(n26485), .ip2(n26484), .ip3(n26483), .ip4(n26482), 
        .op(n26486) );
  not_ab_or_c_or_d U30496 ( .ip1(\LUT[102][10] ), .ip2(n27326), .ip3(n26487), 
        .ip4(n26486), .op(n26491) );
  nand2_1 U30497 ( .ip1(n27370), .ip2(\LUT[100][10] ), .op(n26490) );
  nand2_1 U30498 ( .ip1(n27328), .ip2(\LUT[101][10] ), .op(n26489) );
  nand2_1 U30499 ( .ip1(n27327), .ip2(\LUT[103][10] ), .op(n26488) );
  nand4_1 U30500 ( .ip1(n26491), .ip2(n26490), .ip3(n26489), .ip4(n26488), 
        .op(n26492) );
  not_ab_or_c_or_d U30501 ( .ip1(\LUT[99][10] ), .ip2(n27156), .ip3(n26493), 
        .ip4(n26492), .op(n26494) );
  nor2_1 U30502 ( .ip1(n26494), .ip2(n27371), .op(n26507) );
  nand2_1 U30503 ( .ip1(n27305), .ip2(\LUT[114][10] ), .op(n26498) );
  nand2_1 U30504 ( .ip1(n27298), .ip2(\LUT[117][10] ), .op(n26497) );
  nand2_1 U30505 ( .ip1(n27299), .ip2(\LUT[118][10] ), .op(n26496) );
  nand2_1 U30506 ( .ip1(n27300), .ip2(\LUT[119][10] ), .op(n26495) );
  nand4_1 U30507 ( .ip1(n26498), .ip2(n26497), .ip3(n26496), .ip4(n26495), 
        .op(n26499) );
  or2_1 U30508 ( .ip1(n27297), .ip2(n26499), .op(n26501) );
  or2_1 U30509 ( .ip1(\LUT[116][10] ), .ip2(n26499), .op(n26500) );
  nand2_1 U30510 ( .ip1(n26501), .ip2(n26500), .op(n26505) );
  nand2_1 U30511 ( .ip1(n27172), .ip2(\LUT[111][10] ), .op(n26504) );
  nand2_1 U30512 ( .ip1(n27583), .ip2(\LUT[113][10] ), .op(n26503) );
  nand2_1 U30513 ( .ip1(n27582), .ip2(\LUT[115][10] ), .op(n26502) );
  nand4_1 U30514 ( .ip1(n26505), .ip2(n26504), .ip3(n26503), .ip4(n26502), 
        .op(n26506) );
  not_ab_or_c_or_d U30515 ( .ip1(n27581), .ip2(\LUT[106][10] ), .ip3(n26507), 
        .ip4(n26506), .op(n26625) );
  and2_1 U30516 ( .ip1(n27534), .ip2(\LUT[65][10] ), .op(n26513) );
  nand2_1 U30517 ( .ip1(n27548), .ip2(\LUT[67][10] ), .op(n26511) );
  nand2_1 U30518 ( .ip1(n27536), .ip2(\LUT[70][10] ), .op(n26510) );
  nand2_1 U30519 ( .ip1(n27535), .ip2(\LUT[69][10] ), .op(n26509) );
  nand2_1 U30520 ( .ip1(n27537), .ip2(\LUT[68][10] ), .op(n26508) );
  nand4_1 U30521 ( .ip1(n26511), .ip2(n26510), .ip3(n26509), .ip4(n26508), 
        .op(n26512) );
  not_ab_or_c_or_d U30522 ( .ip1(n27542), .ip2(\LUT[66][10] ), .ip3(n26513), 
        .ip4(n26512), .op(n26517) );
  nand2_1 U30523 ( .ip1(n27547), .ip2(\LUT[64][10] ), .op(n26516) );
  nand2_1 U30524 ( .ip1(n27563), .ip2(\LUT[62][10] ), .op(n26515) );
  nand2_1 U30525 ( .ip1(n27546), .ip2(\LUT[59][10] ), .op(n26514) );
  nand4_1 U30526 ( .ip1(n26517), .ip2(n26516), .ip3(n26515), .ip4(n26514), 
        .op(n26523) );
  nand2_1 U30527 ( .ip1(n27397), .ip2(\LUT[58][10] ), .op(n26521) );
  nand2_1 U30528 ( .ip1(n27556), .ip2(\LUT[63][10] ), .op(n26520) );
  nand2_1 U30529 ( .ip1(n27555), .ip2(\LUT[61][10] ), .op(n26519) );
  nand2_1 U30530 ( .ip1(n27554), .ip2(\LUT[60][10] ), .op(n26518) );
  nand4_1 U30531 ( .ip1(n26521), .ip2(n26520), .ip3(n26519), .ip4(n26518), 
        .op(n26522) );
  not_ab_or_c_or_d U30532 ( .ip1(n27553), .ip2(\LUT[57][10] ), .ip3(n26523), 
        .ip4(n26522), .op(n26524) );
  or2_1 U30533 ( .ip1(n26524), .ip2(n27265), .op(n26602) );
  nand2_1 U30534 ( .ip1(\LUT[27][10] ), .ip2(n27398), .op(n26527) );
  nand2_1 U30535 ( .ip1(n27400), .ip2(\LUT[28][10] ), .op(n26526) );
  nand2_1 U30536 ( .ip1(n27405), .ip2(\LUT[25][10] ), .op(n26525) );
  nand3_1 U30537 ( .ip1(n26527), .ip2(n26526), .ip3(n26525), .op(n26532) );
  nand2_1 U30538 ( .ip1(\LUT[24][10] ), .ip2(n27404), .op(n26530) );
  nand2_1 U30539 ( .ip1(n27399), .ip2(\LUT[26][10] ), .op(n26529) );
  nand2_1 U30540 ( .ip1(n27406), .ip2(\LUT[23][10] ), .op(n26528) );
  nand3_1 U30541 ( .ip1(n26530), .ip2(n26529), .ip3(n26528), .op(n26531) );
  not_ab_or_c_or_d U30542 ( .ip1(n27459), .ip2(\LUT[17][10] ), .ip3(n26532), 
        .ip4(n26531), .op(n26561) );
  nand2_1 U30543 ( .ip1(\LUT[2][10] ), .ip2(n27413), .op(n26534) );
  nand2_1 U30544 ( .ip1(\LUT[3][10] ), .ip2(n27414), .op(n26533) );
  nand2_1 U30545 ( .ip1(n26534), .ip2(n26533), .op(n26550) );
  nand2_1 U30546 ( .ip1(n27428), .ip2(\LUT[6][10] ), .op(n26538) );
  nand2_1 U30547 ( .ip1(n27418), .ip2(\LUT[9][10] ), .op(n26537) );
  nand2_1 U30548 ( .ip1(n27420), .ip2(\LUT[13][10] ), .op(n26536) );
  nand2_1 U30549 ( .ip1(n27419), .ip2(\LUT[14][10] ), .op(n26535) );
  nand4_1 U30550 ( .ip1(n26538), .ip2(n26537), .ip3(n26536), .ip4(n26535), 
        .op(n26544) );
  nand2_1 U30551 ( .ip1(n27426), .ip2(\LUT[8][10] ), .op(n26542) );
  nand2_1 U30552 ( .ip1(n27425), .ip2(\LUT[10][10] ), .op(n26541) );
  nand2_1 U30553 ( .ip1(n27417), .ip2(\LUT[7][10] ), .op(n26540) );
  nand2_1 U30554 ( .ip1(n27427), .ip2(\LUT[12][10] ), .op(n26539) );
  nand4_1 U30555 ( .ip1(n26542), .ip2(n26541), .ip3(n26540), .ip4(n26539), 
        .op(n26543) );
  not_ab_or_c_or_d U30556 ( .ip1(n27435), .ip2(\LUT[11][10] ), .ip3(n26544), 
        .ip4(n26543), .op(n26548) );
  nand2_1 U30557 ( .ip1(n27436), .ip2(\LUT[0][10] ), .op(n26547) );
  nand2_1 U30558 ( .ip1(n27438), .ip2(\LUT[5][10] ), .op(n26546) );
  nand2_1 U30559 ( .ip1(n27437), .ip2(\LUT[4][10] ), .op(n26545) );
  nand4_1 U30560 ( .ip1(n26548), .ip2(n26547), .ip3(n26546), .ip4(n26545), 
        .op(n26549) );
  not_ab_or_c_or_d U30561 ( .ip1(n27445), .ip2(\LUT[1][10] ), .ip3(n26550), 
        .ip4(n26549), .op(n26551) );
  nor2_1 U30562 ( .ip1(n26551), .ip2(n27446), .op(n26557) );
  nand2_1 U30563 ( .ip1(n27451), .ip2(\LUT[16][10] ), .op(n26555) );
  nand2_1 U30564 ( .ip1(n27448), .ip2(\LUT[18][10] ), .op(n26554) );
  nand2_1 U30565 ( .ip1(n27450), .ip2(\LUT[21][10] ), .op(n26553) );
  nand2_1 U30566 ( .ip1(n27449), .ip2(\LUT[20][10] ), .op(n26552) );
  nand4_1 U30567 ( .ip1(n26555), .ip2(n26554), .ip3(n26553), .ip4(n26552), 
        .op(n26556) );
  not_ab_or_c_or_d U30568 ( .ip1(\LUT[15][10] ), .ip2(n27458), .ip3(n26557), 
        .ip4(n26556), .op(n26560) );
  nand2_1 U30569 ( .ip1(n27412), .ip2(\LUT[22][10] ), .op(n26559) );
  nand2_1 U30570 ( .ip1(n27460), .ip2(\LUT[19][10] ), .op(n26558) );
  nand4_1 U30571 ( .ip1(n26561), .ip2(n26560), .ip3(n26559), .ip4(n26558), 
        .op(n26599) );
  nand2_1 U30572 ( .ip1(n27527), .ip2(\LUT[46][10] ), .op(n26565) );
  nand2_1 U30573 ( .ip1(n27498), .ip2(\LUT[48][10] ), .op(n26564) );
  nand2_1 U30574 ( .ip1(n27501), .ip2(\LUT[52][10] ), .op(n26563) );
  nand2_1 U30575 ( .ip1(n27500), .ip2(\LUT[53][10] ), .op(n26562) );
  nand4_1 U30576 ( .ip1(n26565), .ip2(n26564), .ip3(n26563), .ip4(n26562), 
        .op(n26577) );
  and2_1 U30577 ( .ip1(n27518), .ip2(\LUT[44][10] ), .op(n26571) );
  nand2_1 U30578 ( .ip1(n27507), .ip2(\LUT[54][10] ), .op(n26569) );
  nand2_1 U30579 ( .ip1(n27510), .ip2(\LUT[51][10] ), .op(n26568) );
  nand2_1 U30580 ( .ip1(n27509), .ip2(\LUT[56][10] ), .op(n26567) );
  nand2_1 U30581 ( .ip1(n27508), .ip2(\LUT[55][10] ), .op(n26566) );
  nand4_1 U30582 ( .ip1(n26569), .ip2(n26568), .ip3(n26567), .ip4(n26566), 
        .op(n26570) );
  not_ab_or_c_or_d U30583 ( .ip1(\LUT[49][10] ), .ip2(n27499), .ip3(n26571), 
        .ip4(n26570), .op(n26575) );
  nand2_1 U30584 ( .ip1(n27519), .ip2(\LUT[43][10] ), .op(n26574) );
  nand2_1 U30585 ( .ip1(n27506), .ip2(\LUT[45][10] ), .op(n26573) );
  nand2_1 U30586 ( .ip1(n27520), .ip2(\LUT[47][10] ), .op(n26572) );
  nand4_1 U30587 ( .ip1(n26575), .ip2(n26574), .ip3(n26573), .ip4(n26572), 
        .op(n26576) );
  not_ab_or_c_or_d U30588 ( .ip1(n27517), .ip2(\LUT[50][10] ), .ip3(n26577), 
        .ip4(n26576), .op(n26578) );
  nor2_1 U30589 ( .ip1(n26578), .ip2(n27528), .op(n26598) );
  nand2_1 U30590 ( .ip1(\LUT[31][10] ), .ip2(n27465), .op(n26580) );
  nand2_1 U30591 ( .ip1(\LUT[30][10] ), .ip2(n27466), .op(n26579) );
  nand2_1 U30592 ( .ip1(n26580), .ip2(n26579), .op(n26595) );
  nand2_1 U30593 ( .ip1(n27469), .ip2(\LUT[39][10] ), .op(n26584) );
  nand2_1 U30594 ( .ip1(n27470), .ip2(\LUT[38][10] ), .op(n26583) );
  nand2_1 U30595 ( .ip1(n27472), .ip2(\LUT[42][10] ), .op(n26582) );
  nand2_1 U30596 ( .ip1(n27471), .ip2(\LUT[41][10] ), .op(n26581) );
  nand4_1 U30597 ( .ip1(n26584), .ip2(n26583), .ip3(n26582), .ip4(n26581), 
        .op(n26589) );
  nand2_1 U30598 ( .ip1(\LUT[36][10] ), .ip2(n27477), .op(n26587) );
  nand2_1 U30599 ( .ip1(n27488), .ip2(\LUT[33][10] ), .op(n26586) );
  nand2_1 U30600 ( .ip1(n27478), .ip2(\LUT[37][10] ), .op(n26585) );
  nand3_1 U30601 ( .ip1(n26587), .ip2(n26586), .ip3(n26585), .op(n26588) );
  not_ab_or_c_or_d U30602 ( .ip1(n27485), .ip2(\LUT[40][10] ), .ip3(n26589), 
        .ip4(n26588), .op(n26593) );
  nand2_1 U30603 ( .ip1(n27479), .ip2(\LUT[32][10] ), .op(n26592) );
  nand2_1 U30604 ( .ip1(n27487), .ip2(\LUT[35][10] ), .op(n26591) );
  nand2_1 U30605 ( .ip1(n27486), .ip2(\LUT[34][10] ), .op(n26590) );
  nand4_1 U30606 ( .ip1(n26593), .ip2(n26592), .ip3(n26591), .ip4(n26590), 
        .op(n26594) );
  not_ab_or_c_or_d U30607 ( .ip1(n27495), .ip2(\LUT[29][10] ), .ip3(n26595), 
        .ip4(n26594), .op(n26596) );
  nor2_1 U30608 ( .ip1(n26596), .ip2(n27496), .op(n26597) );
  not_ab_or_c_or_d U30609 ( .ip1(n27533), .ip2(n26599), .ip3(n26598), .ip4(
        n26597), .op(n26600) );
  or2_1 U30610 ( .ip1(n26600), .ip2(n27265), .op(n26601) );
  nand2_1 U30611 ( .ip1(n26602), .ip2(n26601), .op(n26616) );
  nand2_1 U30612 ( .ip1(n27391), .ip2(\LUT[75][10] ), .op(n26614) );
  nand2_1 U30613 ( .ip1(n27373), .ip2(\LUT[82][10] ), .op(n26606) );
  nand2_1 U30614 ( .ip1(n27374), .ip2(\LUT[81][10] ), .op(n26605) );
  nand2_1 U30615 ( .ip1(n27376), .ip2(\LUT[83][10] ), .op(n26604) );
  nand2_1 U30616 ( .ip1(n27375), .ip2(\LUT[84][10] ), .op(n26603) );
  nand4_1 U30617 ( .ip1(n26606), .ip2(n26605), .ip3(n26604), .ip4(n26603), 
        .op(n26611) );
  nand2_1 U30618 ( .ip1(\LUT[78][10] ), .ip2(n27381), .op(n26609) );
  nand2_1 U30619 ( .ip1(n27382), .ip2(\LUT[79][10] ), .op(n26608) );
  nand2_1 U30620 ( .ip1(n27383), .ip2(\LUT[77][10] ), .op(n26607) );
  nand3_1 U30621 ( .ip1(n26609), .ip2(n26608), .ip3(n26607), .op(n26610) );
  not_ab_or_c_or_d U30622 ( .ip1(n27389), .ip2(\LUT[80][10] ), .ip3(n26611), 
        .ip4(n26610), .op(n26613) );
  nand2_1 U30623 ( .ip1(n27392), .ip2(\LUT[74][10] ), .op(n26612) );
  nand3_1 U30624 ( .ip1(n26614), .ip2(n26613), .ip3(n26612), .op(n26615) );
  not_ab_or_c_or_d U30625 ( .ip1(n27390), .ip2(\LUT[76][10] ), .ip3(n26616), 
        .ip4(n26615), .op(n26620) );
  nand2_1 U30626 ( .ip1(n27576), .ip2(\LUT[71][10] ), .op(n26619) );
  nand2_1 U30627 ( .ip1(n27570), .ip2(\LUT[72][10] ), .op(n26618) );
  nand2_1 U30628 ( .ip1(n27569), .ip2(\LUT[73][10] ), .op(n26617) );
  nand4_1 U30629 ( .ip1(n26620), .ip2(n26619), .ip3(n26618), .ip4(n26617), 
        .op(n26621) );
  nand2_1 U30630 ( .ip1(n27288), .ip2(n26621), .op(n26624) );
  nand2_1 U30631 ( .ip1(n27289), .ip2(\LUT[112][10] ), .op(n26623) );
  nand2_1 U30632 ( .ip1(n27165), .ip2(\LUT[108][10] ), .op(n26622) );
  nand4_1 U30633 ( .ip1(n26625), .ip2(n26624), .ip3(n26623), .ip4(n26622), 
        .op(n26626) );
  nand2_1 U30634 ( .ip1(n27589), .ip2(n26626), .op(n26628) );
  nand2_1 U30635 ( .ip1(sig_out[10]), .ip2(n27590), .op(n26627) );
  nand2_1 U30636 ( .ip1(n26628), .ip2(n26627), .op(n13455) );
  nand2_1 U30637 ( .ip1(n27333), .ip2(\LUT[95][11] ), .op(n26632) );
  nand2_1 U30638 ( .ip1(n27334), .ip2(\LUT[94][11] ), .op(n26631) );
  nand2_1 U30639 ( .ip1(n27335), .ip2(\LUT[98][11] ), .op(n26630) );
  nand2_1 U30640 ( .ip1(n27336), .ip2(\LUT[97][11] ), .op(n26629) );
  nand4_1 U30641 ( .ip1(n26632), .ip2(n26631), .ip3(n26630), .ip4(n26629), 
        .op(n26637) );
  nand2_1 U30642 ( .ip1(n27341), .ip2(\LUT[93][11] ), .op(n26635) );
  nand2_1 U30643 ( .ip1(n27342), .ip2(\LUT[92][11] ), .op(n26634) );
  nand2_1 U30644 ( .ip1(n27343), .ip2(\LUT[91][11] ), .op(n26633) );
  nand3_1 U30645 ( .ip1(n26635), .ip2(n26634), .ip3(n26633), .op(n26636) );
  not_ab_or_c_or_d U30646 ( .ip1(n27349), .ip2(\LUT[96][11] ), .ip3(n26637), 
        .ip4(n26636), .op(n26641) );
  nand2_1 U30647 ( .ip1(n27350), .ip2(\LUT[89][11] ), .op(n26640) );
  nand2_1 U30648 ( .ip1(n27351), .ip2(\LUT[90][11] ), .op(n26639) );
  nand2_1 U30649 ( .ip1(n27352), .ip2(\LUT[88][11] ), .op(n26638) );
  nand4_1 U30650 ( .ip1(n26641), .ip2(n26640), .ip3(n26639), .ip4(n26638), 
        .op(n26645) );
  nand2_1 U30651 ( .ip1(\LUT[85][11] ), .ip2(n27357), .op(n26643) );
  nand2_1 U30652 ( .ip1(\LUT[86][11] ), .ip2(n27358), .op(n26642) );
  nand2_1 U30653 ( .ip1(n26643), .ip2(n26642), .op(n26644) );
  not_ab_or_c_or_d U30654 ( .ip1(n27363), .ip2(\LUT[87][11] ), .ip3(n26645), 
        .ip4(n26644), .op(n26646) );
  nor2_1 U30655 ( .ip1(n26646), .ip2(n27142), .op(n26660) );
  nand2_1 U30656 ( .ip1(\LUT[110][11] ), .ip2(n27325), .op(n26649) );
  nand2_1 U30657 ( .ip1(n27309), .ip2(\LUT[109][11] ), .op(n26648) );
  nand2_1 U30658 ( .ip1(n27310), .ip2(\LUT[108][11] ), .op(n26647) );
  nand3_1 U30659 ( .ip1(n26649), .ip2(n26648), .ip3(n26647), .op(n26654) );
  nand2_1 U30660 ( .ip1(n27317), .ip2(\LUT[105][11] ), .op(n26652) );
  nand2_1 U30661 ( .ip1(n27318), .ip2(\LUT[107][11] ), .op(n26651) );
  nand2_1 U30662 ( .ip1(n27319), .ip2(\LUT[104][11] ), .op(n26650) );
  nand3_1 U30663 ( .ip1(n26652), .ip2(n26651), .ip3(n26650), .op(n26653) );
  not_ab_or_c_or_d U30664 ( .ip1(n27326), .ip2(\LUT[102][11] ), .ip3(n26654), 
        .ip4(n26653), .op(n26658) );
  nand2_1 U30665 ( .ip1(n27370), .ip2(\LUT[100][11] ), .op(n26657) );
  nand2_1 U30666 ( .ip1(n27328), .ip2(\LUT[101][11] ), .op(n26656) );
  nand2_1 U30667 ( .ip1(n27327), .ip2(\LUT[103][11] ), .op(n26655) );
  nand4_1 U30668 ( .ip1(n26658), .ip2(n26657), .ip3(n26656), .ip4(n26655), 
        .op(n26659) );
  not_ab_or_c_or_d U30669 ( .ip1(\LUT[99][11] ), .ip2(n27156), .ip3(n26660), 
        .ip4(n26659), .op(n26661) );
  nor2_1 U30670 ( .ip1(n26661), .ip2(n27371), .op(n26671) );
  nand2_1 U30671 ( .ip1(n27298), .ip2(\LUT[117][11] ), .op(n26665) );
  nand2_1 U30672 ( .ip1(n27582), .ip2(\LUT[115][11] ), .op(n26664) );
  nand2_1 U30673 ( .ip1(n27300), .ip2(\LUT[119][11] ), .op(n26663) );
  nand2_1 U30674 ( .ip1(n27299), .ip2(\LUT[118][11] ), .op(n26662) );
  and4_1 U30675 ( .ip1(n26665), .ip2(n26664), .ip3(n26663), .ip4(n26662), .op(
        n26669) );
  nand2_1 U30676 ( .ip1(n27289), .ip2(\LUT[112][11] ), .op(n26668) );
  nand2_1 U30677 ( .ip1(n27305), .ip2(\LUT[114][11] ), .op(n26667) );
  nand2_1 U30678 ( .ip1(n27297), .ip2(\LUT[116][11] ), .op(n26666) );
  nand4_1 U30679 ( .ip1(n26669), .ip2(n26668), .ip3(n26667), .ip4(n26666), 
        .op(n26670) );
  not_ab_or_c_or_d U30680 ( .ip1(n27583), .ip2(\LUT[113][11] ), .ip3(n26671), 
        .ip4(n26670), .op(n26791) );
  nand2_1 U30681 ( .ip1(\LUT[27][11] ), .ip2(n27398), .op(n26674) );
  nand2_1 U30682 ( .ip1(n27400), .ip2(\LUT[28][11] ), .op(n26673) );
  nand2_1 U30683 ( .ip1(n27405), .ip2(\LUT[25][11] ), .op(n26672) );
  nand3_1 U30684 ( .ip1(n26674), .ip2(n26673), .ip3(n26672), .op(n26679) );
  nand2_1 U30685 ( .ip1(n27404), .ip2(\LUT[24][11] ), .op(n26677) );
  nand2_1 U30686 ( .ip1(n27406), .ip2(\LUT[23][11] ), .op(n26676) );
  nand2_1 U30687 ( .ip1(n27399), .ip2(\LUT[26][11] ), .op(n26675) );
  nand3_1 U30688 ( .ip1(n26677), .ip2(n26676), .ip3(n26675), .op(n26678) );
  not_ab_or_c_or_d U30689 ( .ip1(n27459), .ip2(\LUT[17][11] ), .ip3(n26679), 
        .ip4(n26678), .op(n26708) );
  nand2_1 U30690 ( .ip1(\LUT[2][11] ), .ip2(n27413), .op(n26681) );
  nand2_1 U30691 ( .ip1(\LUT[3][11] ), .ip2(n27414), .op(n26680) );
  nand2_1 U30692 ( .ip1(n26681), .ip2(n26680), .op(n26697) );
  nand2_1 U30693 ( .ip1(n27428), .ip2(\LUT[6][11] ), .op(n26685) );
  nand2_1 U30694 ( .ip1(n27427), .ip2(\LUT[12][11] ), .op(n26684) );
  nand2_1 U30695 ( .ip1(n27419), .ip2(\LUT[14][11] ), .op(n26683) );
  nand2_1 U30696 ( .ip1(n27420), .ip2(\LUT[13][11] ), .op(n26682) );
  nand4_1 U30697 ( .ip1(n26685), .ip2(n26684), .ip3(n26683), .ip4(n26682), 
        .op(n26691) );
  nand2_1 U30698 ( .ip1(n27417), .ip2(\LUT[7][11] ), .op(n26689) );
  nand2_1 U30699 ( .ip1(n27435), .ip2(\LUT[11][11] ), .op(n26688) );
  nand2_1 U30700 ( .ip1(n27426), .ip2(\LUT[8][11] ), .op(n26687) );
  nand2_1 U30701 ( .ip1(n27425), .ip2(\LUT[10][11] ), .op(n26686) );
  nand4_1 U30702 ( .ip1(n26689), .ip2(n26688), .ip3(n26687), .ip4(n26686), 
        .op(n26690) );
  not_ab_or_c_or_d U30703 ( .ip1(n27418), .ip2(\LUT[9][11] ), .ip3(n26691), 
        .ip4(n26690), .op(n26695) );
  nand2_1 U30704 ( .ip1(n27436), .ip2(\LUT[0][11] ), .op(n26694) );
  nand2_1 U30705 ( .ip1(n27437), .ip2(\LUT[4][11] ), .op(n26693) );
  nand2_1 U30706 ( .ip1(n27438), .ip2(\LUT[5][11] ), .op(n26692) );
  nand4_1 U30707 ( .ip1(n26695), .ip2(n26694), .ip3(n26693), .ip4(n26692), 
        .op(n26696) );
  not_ab_or_c_or_d U30708 ( .ip1(n27445), .ip2(\LUT[1][11] ), .ip3(n26697), 
        .ip4(n26696), .op(n26698) );
  nor2_1 U30709 ( .ip1(n26698), .ip2(n27446), .op(n26704) );
  nand2_1 U30710 ( .ip1(n27451), .ip2(\LUT[16][11] ), .op(n26702) );
  nand2_1 U30711 ( .ip1(n27448), .ip2(\LUT[18][11] ), .op(n26701) );
  nand2_1 U30712 ( .ip1(n27450), .ip2(\LUT[21][11] ), .op(n26700) );
  nand2_1 U30713 ( .ip1(n27449), .ip2(\LUT[20][11] ), .op(n26699) );
  nand4_1 U30714 ( .ip1(n26702), .ip2(n26701), .ip3(n26700), .ip4(n26699), 
        .op(n26703) );
  not_ab_or_c_or_d U30715 ( .ip1(\LUT[15][11] ), .ip2(n27458), .ip3(n26704), 
        .ip4(n26703), .op(n26707) );
  nand2_1 U30716 ( .ip1(n27412), .ip2(\LUT[22][11] ), .op(n26706) );
  nand2_1 U30717 ( .ip1(n27460), .ip2(\LUT[19][11] ), .op(n26705) );
  nand4_1 U30718 ( .ip1(n26708), .ip2(n26707), .ip3(n26706), .ip4(n26705), 
        .op(n26767) );
  nand2_1 U30719 ( .ip1(n27554), .ip2(\LUT[60][11] ), .op(n26712) );
  nand2_1 U30720 ( .ip1(n27397), .ip2(\LUT[58][11] ), .op(n26711) );
  nand2_1 U30721 ( .ip1(n27555), .ip2(\LUT[61][11] ), .op(n26710) );
  nand2_1 U30722 ( .ip1(n27563), .ip2(\LUT[62][11] ), .op(n26709) );
  nand4_1 U30723 ( .ip1(n26712), .ip2(n26711), .ip3(n26710), .ip4(n26709), 
        .op(n26766) );
  nand2_1 U30724 ( .ip1(n27536), .ip2(\LUT[70][11] ), .op(n26716) );
  nand2_1 U30725 ( .ip1(n27535), .ip2(\LUT[69][11] ), .op(n26715) );
  nand2_1 U30726 ( .ip1(n27537), .ip2(\LUT[68][11] ), .op(n26714) );
  nand2_1 U30727 ( .ip1(n27548), .ip2(\LUT[67][11] ), .op(n26713) );
  nand4_1 U30728 ( .ip1(n26716), .ip2(n26715), .ip3(n26714), .ip4(n26713), 
        .op(n26721) );
  nand2_1 U30729 ( .ip1(\LUT[64][11] ), .ip2(n27547), .op(n26719) );
  nand2_1 U30730 ( .ip1(n27542), .ip2(\LUT[66][11] ), .op(n26718) );
  nand2_1 U30731 ( .ip1(n27534), .ip2(\LUT[65][11] ), .op(n26717) );
  nand3_1 U30732 ( .ip1(n26719), .ip2(n26718), .ip3(n26717), .op(n26720) );
  not_ab_or_c_or_d U30733 ( .ip1(n27556), .ip2(\LUT[63][11] ), .ip3(n26721), 
        .ip4(n26720), .op(n26764) );
  nand2_1 U30734 ( .ip1(n27506), .ip2(\LUT[45][11] ), .op(n26725) );
  nand2_1 U30735 ( .ip1(n27500), .ip2(\LUT[53][11] ), .op(n26724) );
  nand2_1 U30736 ( .ip1(n27501), .ip2(\LUT[52][11] ), .op(n26723) );
  nand2_1 U30737 ( .ip1(n27517), .ip2(\LUT[50][11] ), .op(n26722) );
  and4_1 U30738 ( .ip1(n26725), .ip2(n26724), .ip3(n26723), .ip4(n26722), .op(
        n26758) );
  nand2_1 U30739 ( .ip1(\LUT[31][11] ), .ip2(n27465), .op(n26727) );
  nand2_1 U30740 ( .ip1(\LUT[30][11] ), .ip2(n27466), .op(n26726) );
  nand2_1 U30741 ( .ip1(n26727), .ip2(n26726), .op(n26742) );
  nand2_1 U30742 ( .ip1(n27469), .ip2(\LUT[39][11] ), .op(n26731) );
  nand2_1 U30743 ( .ip1(n27470), .ip2(\LUT[38][11] ), .op(n26730) );
  nand2_1 U30744 ( .ip1(n27472), .ip2(\LUT[42][11] ), .op(n26729) );
  nand2_1 U30745 ( .ip1(n27471), .ip2(\LUT[41][11] ), .op(n26728) );
  nand4_1 U30746 ( .ip1(n26731), .ip2(n26730), .ip3(n26729), .ip4(n26728), 
        .op(n26736) );
  nand2_1 U30747 ( .ip1(\LUT[36][11] ), .ip2(n27477), .op(n26734) );
  nand2_1 U30748 ( .ip1(n27478), .ip2(\LUT[37][11] ), .op(n26733) );
  nand2_1 U30749 ( .ip1(n27479), .ip2(\LUT[32][11] ), .op(n26732) );
  nand3_1 U30750 ( .ip1(n26734), .ip2(n26733), .ip3(n26732), .op(n26735) );
  not_ab_or_c_or_d U30751 ( .ip1(n27485), .ip2(\LUT[40][11] ), .ip3(n26736), 
        .ip4(n26735), .op(n26740) );
  nand2_1 U30752 ( .ip1(n27486), .ip2(\LUT[34][11] ), .op(n26739) );
  nand2_1 U30753 ( .ip1(n27488), .ip2(\LUT[33][11] ), .op(n26738) );
  nand2_1 U30754 ( .ip1(n27487), .ip2(\LUT[35][11] ), .op(n26737) );
  nand4_1 U30755 ( .ip1(n26740), .ip2(n26739), .ip3(n26738), .ip4(n26737), 
        .op(n26741) );
  not_ab_or_c_or_d U30756 ( .ip1(n27495), .ip2(\LUT[29][11] ), .ip3(n26742), 
        .ip4(n26741), .op(n26744) );
  nor2_1 U30757 ( .ip1(n26744), .ip2(n26743), .op(n26754) );
  nand2_1 U30758 ( .ip1(n27507), .ip2(\LUT[54][11] ), .op(n26748) );
  nand2_1 U30759 ( .ip1(n27508), .ip2(\LUT[55][11] ), .op(n26747) );
  nand2_1 U30760 ( .ip1(n27509), .ip2(\LUT[56][11] ), .op(n26746) );
  nand2_1 U30761 ( .ip1(n27510), .ip2(\LUT[51][11] ), .op(n26745) );
  and4_1 U30762 ( .ip1(n26748), .ip2(n26747), .ip3(n26746), .ip4(n26745), .op(
        n26752) );
  nand2_1 U30763 ( .ip1(n27520), .ip2(\LUT[47][11] ), .op(n26751) );
  nand2_1 U30764 ( .ip1(n27518), .ip2(\LUT[44][11] ), .op(n26750) );
  nand2_1 U30765 ( .ip1(n27499), .ip2(\LUT[49][11] ), .op(n26749) );
  nand4_1 U30766 ( .ip1(n26752), .ip2(n26751), .ip3(n26750), .ip4(n26749), 
        .op(n26753) );
  not_ab_or_c_or_d U30767 ( .ip1(\LUT[43][11] ), .ip2(n27519), .ip3(n26754), 
        .ip4(n26753), .op(n26757) );
  nand2_1 U30768 ( .ip1(n27498), .ip2(\LUT[48][11] ), .op(n26756) );
  nand2_1 U30769 ( .ip1(n27527), .ip2(\LUT[46][11] ), .op(n26755) );
  nand4_1 U30770 ( .ip1(n26758), .ip2(n26757), .ip3(n26756), .ip4(n26755), 
        .op(n26759) );
  nand2_1 U30771 ( .ip1(n26760), .ip2(n26759), .op(n26763) );
  nand2_1 U30772 ( .ip1(n27553), .ip2(\LUT[57][11] ), .op(n26762) );
  nand2_1 U30773 ( .ip1(n27546), .ip2(\LUT[59][11] ), .op(n26761) );
  nand4_1 U30774 ( .ip1(n26764), .ip2(n26763), .ip3(n26762), .ip4(n26761), 
        .op(n26765) );
  not_ab_or_c_or_d U30775 ( .ip1(n27533), .ip2(n26767), .ip3(n26766), .ip4(
        n26765), .op(n26768) );
  nor2_1 U30776 ( .ip1(n26768), .ip2(n27265), .op(n26782) );
  nand2_1 U30777 ( .ip1(n27391), .ip2(\LUT[75][11] ), .op(n26780) );
  nand2_1 U30778 ( .ip1(n27373), .ip2(\LUT[82][11] ), .op(n26772) );
  nand2_1 U30779 ( .ip1(n27374), .ip2(\LUT[81][11] ), .op(n26771) );
  nand2_1 U30780 ( .ip1(n27375), .ip2(\LUT[84][11] ), .op(n26770) );
  nand2_1 U30781 ( .ip1(n27376), .ip2(\LUT[83][11] ), .op(n26769) );
  nand4_1 U30782 ( .ip1(n26772), .ip2(n26771), .ip3(n26770), .ip4(n26769), 
        .op(n26777) );
  nand2_1 U30783 ( .ip1(\LUT[78][11] ), .ip2(n27381), .op(n26775) );
  nand2_1 U30784 ( .ip1(n27382), .ip2(\LUT[79][11] ), .op(n26774) );
  nand2_1 U30785 ( .ip1(n27383), .ip2(\LUT[77][11] ), .op(n26773) );
  nand3_1 U30786 ( .ip1(n26775), .ip2(n26774), .ip3(n26773), .op(n26776) );
  not_ab_or_c_or_d U30787 ( .ip1(n27389), .ip2(\LUT[80][11] ), .ip3(n26777), 
        .ip4(n26776), .op(n26779) );
  nand2_1 U30788 ( .ip1(n27392), .ip2(\LUT[74][11] ), .op(n26778) );
  nand3_1 U30789 ( .ip1(n26780), .ip2(n26779), .ip3(n26778), .op(n26781) );
  not_ab_or_c_or_d U30790 ( .ip1(n27390), .ip2(\LUT[76][11] ), .ip3(n26782), 
        .ip4(n26781), .op(n26786) );
  nand2_1 U30791 ( .ip1(n27576), .ip2(\LUT[71][11] ), .op(n26785) );
  nand2_1 U30792 ( .ip1(n27570), .ip2(\LUT[72][11] ), .op(n26784) );
  nand2_1 U30793 ( .ip1(n27569), .ip2(\LUT[73][11] ), .op(n26783) );
  nand4_1 U30794 ( .ip1(n26786), .ip2(n26785), .ip3(n26784), .ip4(n26783), 
        .op(n26787) );
  nand2_1 U30795 ( .ip1(n27288), .ip2(n26787), .op(n26790) );
  nand2_1 U30796 ( .ip1(n27581), .ip2(\LUT[106][11] ), .op(n26789) );
  nand2_1 U30797 ( .ip1(n27172), .ip2(\LUT[111][11] ), .op(n26788) );
  nand4_1 U30798 ( .ip1(n26791), .ip2(n26790), .ip3(n26789), .ip4(n26788), 
        .op(n26792) );
  nand2_1 U30799 ( .ip1(n27589), .ip2(n26792), .op(n26794) );
  nand2_1 U30800 ( .ip1(sig_out[11]), .ip2(n27590), .op(n26793) );
  nand2_1 U30801 ( .ip1(n26794), .ip2(n26793), .op(n13454) );
  nand2_1 U30802 ( .ip1(n27333), .ip2(\LUT[95][12] ), .op(n26798) );
  nand2_1 U30803 ( .ip1(n27334), .ip2(\LUT[94][12] ), .op(n26797) );
  nand2_1 U30804 ( .ip1(n27335), .ip2(\LUT[98][12] ), .op(n26796) );
  nand2_1 U30805 ( .ip1(n27336), .ip2(\LUT[97][12] ), .op(n26795) );
  nand4_1 U30806 ( .ip1(n26798), .ip2(n26797), .ip3(n26796), .ip4(n26795), 
        .op(n26803) );
  nand2_1 U30807 ( .ip1(n27341), .ip2(\LUT[93][12] ), .op(n26801) );
  nand2_1 U30808 ( .ip1(n27342), .ip2(\LUT[92][12] ), .op(n26800) );
  nand2_1 U30809 ( .ip1(n27343), .ip2(\LUT[91][12] ), .op(n26799) );
  nand3_1 U30810 ( .ip1(n26801), .ip2(n26800), .ip3(n26799), .op(n26802) );
  not_ab_or_c_or_d U30811 ( .ip1(n27349), .ip2(\LUT[96][12] ), .ip3(n26803), 
        .ip4(n26802), .op(n26807) );
  nand2_1 U30812 ( .ip1(n27350), .ip2(\LUT[89][12] ), .op(n26806) );
  nand2_1 U30813 ( .ip1(n27351), .ip2(\LUT[90][12] ), .op(n26805) );
  nand2_1 U30814 ( .ip1(n27352), .ip2(\LUT[88][12] ), .op(n26804) );
  nand4_1 U30815 ( .ip1(n26807), .ip2(n26806), .ip3(n26805), .ip4(n26804), 
        .op(n26811) );
  nand2_1 U30816 ( .ip1(\LUT[85][12] ), .ip2(n27357), .op(n26809) );
  nand2_1 U30817 ( .ip1(\LUT[86][12] ), .ip2(n27358), .op(n26808) );
  nand2_1 U30818 ( .ip1(n26809), .ip2(n26808), .op(n26810) );
  not_ab_or_c_or_d U30819 ( .ip1(n27363), .ip2(\LUT[87][12] ), .ip3(n26811), 
        .ip4(n26810), .op(n26812) );
  nor2_1 U30820 ( .ip1(n26812), .ip2(n27142), .op(n26824) );
  and2_1 U30821 ( .ip1(n27317), .ip2(\LUT[105][12] ), .op(n26818) );
  nand2_1 U30822 ( .ip1(n27318), .ip2(\LUT[107][12] ), .op(n26816) );
  nand2_1 U30823 ( .ip1(n27319), .ip2(\LUT[104][12] ), .op(n26815) );
  nand2_1 U30824 ( .ip1(n27325), .ip2(\LUT[110][12] ), .op(n26814) );
  nand2_1 U30825 ( .ip1(n27309), .ip2(\LUT[109][12] ), .op(n26813) );
  nand4_1 U30826 ( .ip1(n26816), .ip2(n26815), .ip3(n26814), .ip4(n26813), 
        .op(n26817) );
  not_ab_or_c_or_d U30827 ( .ip1(\LUT[102][12] ), .ip2(n27326), .ip3(n26818), 
        .ip4(n26817), .op(n26822) );
  nand2_1 U30828 ( .ip1(n27370), .ip2(\LUT[100][12] ), .op(n26821) );
  nand2_1 U30829 ( .ip1(n27328), .ip2(\LUT[101][12] ), .op(n26820) );
  nand2_1 U30830 ( .ip1(n27327), .ip2(\LUT[103][12] ), .op(n26819) );
  nand4_1 U30831 ( .ip1(n26822), .ip2(n26821), .ip3(n26820), .ip4(n26819), 
        .op(n26823) );
  not_ab_or_c_or_d U30832 ( .ip1(\LUT[99][12] ), .ip2(n27156), .ip3(n26824), 
        .ip4(n26823), .op(n26825) );
  nor2_1 U30833 ( .ip1(n26825), .ip2(n27371), .op(n26838) );
  nand2_1 U30834 ( .ip1(n27582), .ip2(\LUT[115][12] ), .op(n26829) );
  nand2_1 U30835 ( .ip1(n27298), .ip2(\LUT[117][12] ), .op(n26828) );
  nand2_1 U30836 ( .ip1(n27299), .ip2(\LUT[118][12] ), .op(n26827) );
  nand2_1 U30837 ( .ip1(n27300), .ip2(\LUT[119][12] ), .op(n26826) );
  nand4_1 U30838 ( .ip1(n26829), .ip2(n26828), .ip3(n26827), .ip4(n26826), 
        .op(n26830) );
  or2_1 U30839 ( .ip1(n27297), .ip2(n26830), .op(n26832) );
  or2_1 U30840 ( .ip1(\LUT[116][12] ), .ip2(n26830), .op(n26831) );
  nand2_1 U30841 ( .ip1(n26832), .ip2(n26831), .op(n26836) );
  nand2_1 U30842 ( .ip1(n27165), .ip2(\LUT[108][12] ), .op(n26835) );
  nand2_1 U30843 ( .ip1(n27289), .ip2(\LUT[112][12] ), .op(n26834) );
  nand2_1 U30844 ( .ip1(n27305), .ip2(\LUT[114][12] ), .op(n26833) );
  nand4_1 U30845 ( .ip1(n26836), .ip2(n26835), .ip3(n26834), .ip4(n26833), 
        .op(n26837) );
  not_ab_or_c_or_d U30846 ( .ip1(n27583), .ip2(\LUT[113][12] ), .ip3(n26838), 
        .ip4(n26837), .op(n26956) );
  and2_1 U30847 ( .ip1(n27534), .ip2(\LUT[65][12] ), .op(n26844) );
  nand2_1 U30848 ( .ip1(n27548), .ip2(\LUT[67][12] ), .op(n26842) );
  nand2_1 U30849 ( .ip1(n27537), .ip2(\LUT[68][12] ), .op(n26841) );
  nand2_1 U30850 ( .ip1(n27535), .ip2(\LUT[69][12] ), .op(n26840) );
  nand2_1 U30851 ( .ip1(n27536), .ip2(\LUT[70][12] ), .op(n26839) );
  nand4_1 U30852 ( .ip1(n26842), .ip2(n26841), .ip3(n26840), .ip4(n26839), 
        .op(n26843) );
  not_ab_or_c_or_d U30853 ( .ip1(n27542), .ip2(\LUT[66][12] ), .ip3(n26844), 
        .ip4(n26843), .op(n26848) );
  nand2_1 U30854 ( .ip1(n27546), .ip2(\LUT[59][12] ), .op(n26847) );
  nand2_1 U30855 ( .ip1(n27547), .ip2(\LUT[64][12] ), .op(n26846) );
  nand2_1 U30856 ( .ip1(n27555), .ip2(\LUT[61][12] ), .op(n26845) );
  nand4_1 U30857 ( .ip1(n26848), .ip2(n26847), .ip3(n26846), .ip4(n26845), 
        .op(n26854) );
  nand2_1 U30858 ( .ip1(n27553), .ip2(\LUT[57][12] ), .op(n26852) );
  nand2_1 U30859 ( .ip1(n27554), .ip2(\LUT[60][12] ), .op(n26851) );
  nand2_1 U30860 ( .ip1(n27563), .ip2(\LUT[62][12] ), .op(n26850) );
  nand2_1 U30861 ( .ip1(n27556), .ip2(\LUT[63][12] ), .op(n26849) );
  nand4_1 U30862 ( .ip1(n26852), .ip2(n26851), .ip3(n26850), .ip4(n26849), 
        .op(n26853) );
  not_ab_or_c_or_d U30863 ( .ip1(n27397), .ip2(\LUT[58][12] ), .ip3(n26854), 
        .ip4(n26853), .op(n26855) );
  or2_1 U30864 ( .ip1(n26855), .ip2(n27265), .op(n26933) );
  nand2_1 U30865 ( .ip1(\LUT[27][12] ), .ip2(n27398), .op(n26858) );
  nand2_1 U30866 ( .ip1(n27399), .ip2(\LUT[26][12] ), .op(n26857) );
  nand2_1 U30867 ( .ip1(n27400), .ip2(\LUT[28][12] ), .op(n26856) );
  nand3_1 U30868 ( .ip1(n26858), .ip2(n26857), .ip3(n26856), .op(n26863) );
  nand2_1 U30869 ( .ip1(n27404), .ip2(\LUT[24][12] ), .op(n26861) );
  nand2_1 U30870 ( .ip1(n27405), .ip2(\LUT[25][12] ), .op(n26860) );
  nand2_1 U30871 ( .ip1(n27406), .ip2(\LUT[23][12] ), .op(n26859) );
  nand3_1 U30872 ( .ip1(n26861), .ip2(n26860), .ip3(n26859), .op(n26862) );
  not_ab_or_c_or_d U30873 ( .ip1(n27412), .ip2(\LUT[22][12] ), .ip3(n26863), 
        .ip4(n26862), .op(n26892) );
  nand2_1 U30874 ( .ip1(\LUT[2][12] ), .ip2(n27413), .op(n26865) );
  nand2_1 U30875 ( .ip1(\LUT[3][12] ), .ip2(n27414), .op(n26864) );
  nand2_1 U30876 ( .ip1(n26865), .ip2(n26864), .op(n26881) );
  nand2_1 U30877 ( .ip1(n27428), .ip2(\LUT[6][12] ), .op(n26869) );
  nand2_1 U30878 ( .ip1(n27418), .ip2(\LUT[9][12] ), .op(n26868) );
  nand2_1 U30879 ( .ip1(n27419), .ip2(\LUT[14][12] ), .op(n26867) );
  nand2_1 U30880 ( .ip1(n27420), .ip2(\LUT[13][12] ), .op(n26866) );
  nand4_1 U30881 ( .ip1(n26869), .ip2(n26868), .ip3(n26867), .ip4(n26866), 
        .op(n26875) );
  nand2_1 U30882 ( .ip1(n27425), .ip2(\LUT[10][12] ), .op(n26873) );
  nand2_1 U30883 ( .ip1(n27417), .ip2(\LUT[7][12] ), .op(n26872) );
  nand2_1 U30884 ( .ip1(n27427), .ip2(\LUT[12][12] ), .op(n26871) );
  nand2_1 U30885 ( .ip1(n27426), .ip2(\LUT[8][12] ), .op(n26870) );
  nand4_1 U30886 ( .ip1(n26873), .ip2(n26872), .ip3(n26871), .ip4(n26870), 
        .op(n26874) );
  not_ab_or_c_or_d U30887 ( .ip1(n27435), .ip2(\LUT[11][12] ), .ip3(n26875), 
        .ip4(n26874), .op(n26879) );
  nand2_1 U30888 ( .ip1(n27436), .ip2(\LUT[0][12] ), .op(n26878) );
  nand2_1 U30889 ( .ip1(n27437), .ip2(\LUT[4][12] ), .op(n26877) );
  nand2_1 U30890 ( .ip1(n27438), .ip2(\LUT[5][12] ), .op(n26876) );
  nand4_1 U30891 ( .ip1(n26879), .ip2(n26878), .ip3(n26877), .ip4(n26876), 
        .op(n26880) );
  not_ab_or_c_or_d U30892 ( .ip1(n27445), .ip2(\LUT[1][12] ), .ip3(n26881), 
        .ip4(n26880), .op(n26882) );
  nor2_1 U30893 ( .ip1(n26882), .ip2(n27446), .op(n26888) );
  nand2_1 U30894 ( .ip1(n27448), .ip2(\LUT[18][12] ), .op(n26886) );
  nand2_1 U30895 ( .ip1(n27450), .ip2(\LUT[21][12] ), .op(n26885) );
  nand2_1 U30896 ( .ip1(n27449), .ip2(\LUT[20][12] ), .op(n26884) );
  nand2_1 U30897 ( .ip1(n27451), .ip2(\LUT[16][12] ), .op(n26883) );
  nand4_1 U30898 ( .ip1(n26886), .ip2(n26885), .ip3(n26884), .ip4(n26883), 
        .op(n26887) );
  not_ab_or_c_or_d U30899 ( .ip1(\LUT[15][12] ), .ip2(n27458), .ip3(n26888), 
        .ip4(n26887), .op(n26891) );
  nand2_1 U30900 ( .ip1(n27459), .ip2(\LUT[17][12] ), .op(n26890) );
  nand2_1 U30901 ( .ip1(n27460), .ip2(\LUT[19][12] ), .op(n26889) );
  nand4_1 U30902 ( .ip1(n26892), .ip2(n26891), .ip3(n26890), .ip4(n26889), 
        .op(n26930) );
  nand2_1 U30903 ( .ip1(n27498), .ip2(\LUT[48][12] ), .op(n26896) );
  nand2_1 U30904 ( .ip1(n27499), .ip2(\LUT[49][12] ), .op(n26895) );
  nand2_1 U30905 ( .ip1(n27500), .ip2(\LUT[53][12] ), .op(n26894) );
  nand2_1 U30906 ( .ip1(n27501), .ip2(\LUT[52][12] ), .op(n26893) );
  nand4_1 U30907 ( .ip1(n26896), .ip2(n26895), .ip3(n26894), .ip4(n26893), 
        .op(n26908) );
  and2_1 U30908 ( .ip1(n27518), .ip2(\LUT[44][12] ), .op(n26902) );
  nand2_1 U30909 ( .ip1(n27507), .ip2(\LUT[54][12] ), .op(n26900) );
  nand2_1 U30910 ( .ip1(n27509), .ip2(\LUT[56][12] ), .op(n26899) );
  nand2_1 U30911 ( .ip1(n27508), .ip2(\LUT[55][12] ), .op(n26898) );
  nand2_1 U30912 ( .ip1(n27510), .ip2(\LUT[51][12] ), .op(n26897) );
  nand4_1 U30913 ( .ip1(n26900), .ip2(n26899), .ip3(n26898), .ip4(n26897), 
        .op(n26901) );
  not_ab_or_c_or_d U30914 ( .ip1(n27517), .ip2(\LUT[50][12] ), .ip3(n26902), 
        .ip4(n26901), .op(n26906) );
  nand2_1 U30915 ( .ip1(n27506), .ip2(\LUT[45][12] ), .op(n26905) );
  nand2_1 U30916 ( .ip1(n27519), .ip2(\LUT[43][12] ), .op(n26904) );
  nand2_1 U30917 ( .ip1(n27520), .ip2(\LUT[47][12] ), .op(n26903) );
  nand4_1 U30918 ( .ip1(n26906), .ip2(n26905), .ip3(n26904), .ip4(n26903), 
        .op(n26907) );
  not_ab_or_c_or_d U30919 ( .ip1(n27527), .ip2(\LUT[46][12] ), .ip3(n26908), 
        .ip4(n26907), .op(n26909) );
  nor2_1 U30920 ( .ip1(n26909), .ip2(n27528), .op(n26929) );
  nand2_1 U30921 ( .ip1(\LUT[31][12] ), .ip2(n27465), .op(n26911) );
  nand2_1 U30922 ( .ip1(\LUT[30][12] ), .ip2(n27466), .op(n26910) );
  nand2_1 U30923 ( .ip1(n26911), .ip2(n26910), .op(n26926) );
  nand2_1 U30924 ( .ip1(n27469), .ip2(\LUT[39][12] ), .op(n26915) );
  nand2_1 U30925 ( .ip1(n27470), .ip2(\LUT[38][12] ), .op(n26914) );
  nand2_1 U30926 ( .ip1(n27471), .ip2(\LUT[41][12] ), .op(n26913) );
  nand2_1 U30927 ( .ip1(n27472), .ip2(\LUT[42][12] ), .op(n26912) );
  nand4_1 U30928 ( .ip1(n26915), .ip2(n26914), .ip3(n26913), .ip4(n26912), 
        .op(n26920) );
  nand2_1 U30929 ( .ip1(\LUT[36][12] ), .ip2(n27477), .op(n26918) );
  nand2_1 U30930 ( .ip1(n27478), .ip2(\LUT[37][12] ), .op(n26917) );
  nand2_1 U30931 ( .ip1(n27479), .ip2(\LUT[32][12] ), .op(n26916) );
  nand3_1 U30932 ( .ip1(n26918), .ip2(n26917), .ip3(n26916), .op(n26919) );
  not_ab_or_c_or_d U30933 ( .ip1(n27485), .ip2(\LUT[40][12] ), .ip3(n26920), 
        .ip4(n26919), .op(n26924) );
  nand2_1 U30934 ( .ip1(n27486), .ip2(\LUT[34][12] ), .op(n26923) );
  nand2_1 U30935 ( .ip1(n27488), .ip2(\LUT[33][12] ), .op(n26922) );
  nand2_1 U30936 ( .ip1(n27487), .ip2(\LUT[35][12] ), .op(n26921) );
  nand4_1 U30937 ( .ip1(n26924), .ip2(n26923), .ip3(n26922), .ip4(n26921), 
        .op(n26925) );
  not_ab_or_c_or_d U30938 ( .ip1(n27495), .ip2(\LUT[29][12] ), .ip3(n26926), 
        .ip4(n26925), .op(n26927) );
  nor2_1 U30939 ( .ip1(n26927), .ip2(n27496), .op(n26928) );
  not_ab_or_c_or_d U30940 ( .ip1(n27533), .ip2(n26930), .ip3(n26929), .ip4(
        n26928), .op(n26931) );
  or2_1 U30941 ( .ip1(n26931), .ip2(n27265), .op(n26932) );
  nand2_1 U30942 ( .ip1(n26933), .ip2(n26932), .op(n26947) );
  nand2_1 U30943 ( .ip1(n27391), .ip2(\LUT[75][12] ), .op(n26945) );
  nand2_1 U30944 ( .ip1(n27373), .ip2(\LUT[82][12] ), .op(n26937) );
  nand2_1 U30945 ( .ip1(n27374), .ip2(\LUT[81][12] ), .op(n26936) );
  nand2_1 U30946 ( .ip1(n27375), .ip2(\LUT[84][12] ), .op(n26935) );
  nand2_1 U30947 ( .ip1(n27376), .ip2(\LUT[83][12] ), .op(n26934) );
  nand4_1 U30948 ( .ip1(n26937), .ip2(n26936), .ip3(n26935), .ip4(n26934), 
        .op(n26942) );
  nand2_1 U30949 ( .ip1(n27381), .ip2(\LUT[78][12] ), .op(n26940) );
  nand2_1 U30950 ( .ip1(n27382), .ip2(\LUT[79][12] ), .op(n26939) );
  nand2_1 U30951 ( .ip1(n27383), .ip2(\LUT[77][12] ), .op(n26938) );
  nand3_1 U30952 ( .ip1(n26940), .ip2(n26939), .ip3(n26938), .op(n26941) );
  not_ab_or_c_or_d U30953 ( .ip1(n27389), .ip2(\LUT[80][12] ), .ip3(n26942), 
        .ip4(n26941), .op(n26944) );
  nand2_1 U30954 ( .ip1(n27392), .ip2(\LUT[74][12] ), .op(n26943) );
  nand3_1 U30955 ( .ip1(n26945), .ip2(n26944), .ip3(n26943), .op(n26946) );
  not_ab_or_c_or_d U30956 ( .ip1(n27390), .ip2(\LUT[76][12] ), .ip3(n26947), 
        .ip4(n26946), .op(n26951) );
  nand2_1 U30957 ( .ip1(n27576), .ip2(\LUT[71][12] ), .op(n26950) );
  nand2_1 U30958 ( .ip1(n27569), .ip2(\LUT[73][12] ), .op(n26949) );
  nand2_1 U30959 ( .ip1(n27570), .ip2(\LUT[72][12] ), .op(n26948) );
  nand4_1 U30960 ( .ip1(n26951), .ip2(n26950), .ip3(n26949), .ip4(n26948), 
        .op(n26952) );
  nand2_1 U30961 ( .ip1(n27288), .ip2(n26952), .op(n26955) );
  nand2_1 U30962 ( .ip1(n27581), .ip2(\LUT[106][12] ), .op(n26954) );
  nand2_1 U30963 ( .ip1(n27172), .ip2(\LUT[111][12] ), .op(n26953) );
  nand4_1 U30964 ( .ip1(n26956), .ip2(n26955), .ip3(n26954), .ip4(n26953), 
        .op(n26957) );
  nand2_1 U30965 ( .ip1(n27589), .ip2(n26957), .op(n26959) );
  nand2_1 U30966 ( .ip1(sig_out[12]), .ip2(n27590), .op(n26958) );
  nand2_1 U30967 ( .ip1(n26959), .ip2(n26958), .op(n13453) );
  nand2_1 U30968 ( .ip1(n27333), .ip2(\LUT[95][13] ), .op(n26963) );
  nand2_1 U30969 ( .ip1(n27334), .ip2(\LUT[94][13] ), .op(n26962) );
  nand2_1 U30970 ( .ip1(n27336), .ip2(\LUT[97][13] ), .op(n26961) );
  nand2_1 U30971 ( .ip1(n27335), .ip2(\LUT[98][13] ), .op(n26960) );
  nand4_1 U30972 ( .ip1(n26963), .ip2(n26962), .ip3(n26961), .ip4(n26960), 
        .op(n26968) );
  nand2_1 U30973 ( .ip1(n27341), .ip2(\LUT[93][13] ), .op(n26966) );
  nand2_1 U30974 ( .ip1(n27342), .ip2(\LUT[92][13] ), .op(n26965) );
  nand2_1 U30975 ( .ip1(n27343), .ip2(\LUT[91][13] ), .op(n26964) );
  nand3_1 U30976 ( .ip1(n26966), .ip2(n26965), .ip3(n26964), .op(n26967) );
  not_ab_or_c_or_d U30977 ( .ip1(n27349), .ip2(\LUT[96][13] ), .ip3(n26968), 
        .ip4(n26967), .op(n26972) );
  nand2_1 U30978 ( .ip1(n27350), .ip2(\LUT[89][13] ), .op(n26971) );
  nand2_1 U30979 ( .ip1(n27351), .ip2(\LUT[90][13] ), .op(n26970) );
  nand2_1 U30980 ( .ip1(n27352), .ip2(\LUT[88][13] ), .op(n26969) );
  nand4_1 U30981 ( .ip1(n26972), .ip2(n26971), .ip3(n26970), .ip4(n26969), 
        .op(n26976) );
  nand2_1 U30982 ( .ip1(\LUT[85][13] ), .ip2(n27357), .op(n26974) );
  nand2_1 U30983 ( .ip1(\LUT[86][13] ), .ip2(n27358), .op(n26973) );
  nand2_1 U30984 ( .ip1(n26974), .ip2(n26973), .op(n26975) );
  not_ab_or_c_or_d U30985 ( .ip1(n27363), .ip2(\LUT[87][13] ), .ip3(n26976), 
        .ip4(n26975), .op(n26977) );
  nor2_1 U30986 ( .ip1(n26977), .ip2(n27142), .op(n26989) );
  and2_1 U30987 ( .ip1(n27317), .ip2(\LUT[105][13] ), .op(n26983) );
  nand2_1 U30988 ( .ip1(n27318), .ip2(\LUT[107][13] ), .op(n26981) );
  nand2_1 U30989 ( .ip1(n27319), .ip2(\LUT[104][13] ), .op(n26980) );
  nand2_1 U30990 ( .ip1(n27309), .ip2(\LUT[109][13] ), .op(n26979) );
  nand2_1 U30991 ( .ip1(n27325), .ip2(\LUT[110][13] ), .op(n26978) );
  nand4_1 U30992 ( .ip1(n26981), .ip2(n26980), .ip3(n26979), .ip4(n26978), 
        .op(n26982) );
  not_ab_or_c_or_d U30993 ( .ip1(\LUT[102][13] ), .ip2(n27326), .ip3(n26983), 
        .ip4(n26982), .op(n26987) );
  nand2_1 U30994 ( .ip1(n27370), .ip2(\LUT[100][13] ), .op(n26986) );
  nand2_1 U30995 ( .ip1(n27328), .ip2(\LUT[101][13] ), .op(n26985) );
  nand2_1 U30996 ( .ip1(n27327), .ip2(\LUT[103][13] ), .op(n26984) );
  nand4_1 U30997 ( .ip1(n26987), .ip2(n26986), .ip3(n26985), .ip4(n26984), 
        .op(n26988) );
  not_ab_or_c_or_d U30998 ( .ip1(\LUT[99][13] ), .ip2(n27156), .ip3(n26989), 
        .ip4(n26988), .op(n26990) );
  nor2_1 U30999 ( .ip1(n26990), .ip2(n27371), .op(n27003) );
  nand2_1 U31000 ( .ip1(n27582), .ip2(\LUT[115][13] ), .op(n26994) );
  nand2_1 U31001 ( .ip1(n27298), .ip2(\LUT[117][13] ), .op(n26993) );
  nand2_1 U31002 ( .ip1(n27299), .ip2(\LUT[118][13] ), .op(n26992) );
  nand2_1 U31003 ( .ip1(n27300), .ip2(\LUT[119][13] ), .op(n26991) );
  nand4_1 U31004 ( .ip1(n26994), .ip2(n26993), .ip3(n26992), .ip4(n26991), 
        .op(n26995) );
  or2_1 U31005 ( .ip1(n27297), .ip2(n26995), .op(n26997) );
  or2_1 U31006 ( .ip1(\LUT[116][13] ), .ip2(n26995), .op(n26996) );
  nand2_1 U31007 ( .ip1(n26997), .ip2(n26996), .op(n27001) );
  nand2_1 U31008 ( .ip1(n27583), .ip2(\LUT[113][13] ), .op(n27000) );
  nand2_1 U31009 ( .ip1(n27165), .ip2(\LUT[108][13] ), .op(n26999) );
  nand2_1 U31010 ( .ip1(n27305), .ip2(\LUT[114][13] ), .op(n26998) );
  nand4_1 U31011 ( .ip1(n27001), .ip2(n27000), .ip3(n26999), .ip4(n26998), 
        .op(n27002) );
  not_ab_or_c_or_d U31012 ( .ip1(n27581), .ip2(\LUT[106][13] ), .ip3(n27003), 
        .ip4(n27002), .op(n27121) );
  and2_1 U31013 ( .ip1(n27548), .ip2(\LUT[67][13] ), .op(n27009) );
  nand2_1 U31014 ( .ip1(n27534), .ip2(\LUT[65][13] ), .op(n27007) );
  nand2_1 U31015 ( .ip1(n27535), .ip2(\LUT[69][13] ), .op(n27006) );
  nand2_1 U31016 ( .ip1(n27536), .ip2(\LUT[70][13] ), .op(n27005) );
  nand2_1 U31017 ( .ip1(n27537), .ip2(\LUT[68][13] ), .op(n27004) );
  nand4_1 U31018 ( .ip1(n27007), .ip2(n27006), .ip3(n27005), .ip4(n27004), 
        .op(n27008) );
  not_ab_or_c_or_d U31019 ( .ip1(n27542), .ip2(\LUT[66][13] ), .ip3(n27009), 
        .ip4(n27008), .op(n27013) );
  nand2_1 U31020 ( .ip1(n27546), .ip2(\LUT[59][13] ), .op(n27012) );
  nand2_1 U31021 ( .ip1(n27547), .ip2(\LUT[64][13] ), .op(n27011) );
  nand2_1 U31022 ( .ip1(n27555), .ip2(\LUT[61][13] ), .op(n27010) );
  nand4_1 U31023 ( .ip1(n27013), .ip2(n27012), .ip3(n27011), .ip4(n27010), 
        .op(n27019) );
  nand2_1 U31024 ( .ip1(n27553), .ip2(\LUT[57][13] ), .op(n27017) );
  nand2_1 U31025 ( .ip1(n27556), .ip2(\LUT[63][13] ), .op(n27016) );
  nand2_1 U31026 ( .ip1(n27554), .ip2(\LUT[60][13] ), .op(n27015) );
  nand2_1 U31027 ( .ip1(n27563), .ip2(\LUT[62][13] ), .op(n27014) );
  nand4_1 U31028 ( .ip1(n27017), .ip2(n27016), .ip3(n27015), .ip4(n27014), 
        .op(n27018) );
  not_ab_or_c_or_d U31029 ( .ip1(n27397), .ip2(\LUT[58][13] ), .ip3(n27019), 
        .ip4(n27018), .op(n27020) );
  or2_1 U31030 ( .ip1(n27020), .ip2(n27265), .op(n27098) );
  nand2_1 U31031 ( .ip1(\LUT[27][13] ), .ip2(n27398), .op(n27023) );
  nand2_1 U31032 ( .ip1(n27399), .ip2(\LUT[26][13] ), .op(n27022) );
  nand2_1 U31033 ( .ip1(n27400), .ip2(\LUT[28][13] ), .op(n27021) );
  nand3_1 U31034 ( .ip1(n27023), .ip2(n27022), .ip3(n27021), .op(n27028) );
  nand2_1 U31035 ( .ip1(n27404), .ip2(\LUT[24][13] ), .op(n27026) );
  nand2_1 U31036 ( .ip1(n27405), .ip2(\LUT[25][13] ), .op(n27025) );
  nand2_1 U31037 ( .ip1(n27406), .ip2(\LUT[23][13] ), .op(n27024) );
  nand3_1 U31038 ( .ip1(n27026), .ip2(n27025), .ip3(n27024), .op(n27027) );
  not_ab_or_c_or_d U31039 ( .ip1(n27412), .ip2(\LUT[22][13] ), .ip3(n27028), 
        .ip4(n27027), .op(n27057) );
  nand2_1 U31040 ( .ip1(\LUT[2][13] ), .ip2(n27413), .op(n27030) );
  nand2_1 U31041 ( .ip1(\LUT[3][13] ), .ip2(n27414), .op(n27029) );
  nand2_1 U31042 ( .ip1(n27030), .ip2(n27029), .op(n27046) );
  nand2_1 U31043 ( .ip1(n27418), .ip2(\LUT[9][13] ), .op(n27034) );
  nand2_1 U31044 ( .ip1(n27417), .ip2(\LUT[7][13] ), .op(n27033) );
  nand2_1 U31045 ( .ip1(n27419), .ip2(\LUT[14][13] ), .op(n27032) );
  nand2_1 U31046 ( .ip1(n27420), .ip2(\LUT[13][13] ), .op(n27031) );
  nand4_1 U31047 ( .ip1(n27034), .ip2(n27033), .ip3(n27032), .ip4(n27031), 
        .op(n27040) );
  nand2_1 U31048 ( .ip1(n27427), .ip2(\LUT[12][13] ), .op(n27038) );
  nand2_1 U31049 ( .ip1(n27428), .ip2(\LUT[6][13] ), .op(n27037) );
  nand2_1 U31050 ( .ip1(n27426), .ip2(\LUT[8][13] ), .op(n27036) );
  nand2_1 U31051 ( .ip1(n27425), .ip2(\LUT[10][13] ), .op(n27035) );
  nand4_1 U31052 ( .ip1(n27038), .ip2(n27037), .ip3(n27036), .ip4(n27035), 
        .op(n27039) );
  not_ab_or_c_or_d U31053 ( .ip1(n27435), .ip2(\LUT[11][13] ), .ip3(n27040), 
        .ip4(n27039), .op(n27044) );
  nand2_1 U31054 ( .ip1(n27445), .ip2(\LUT[1][13] ), .op(n27043) );
  nand2_1 U31055 ( .ip1(n27437), .ip2(\LUT[4][13] ), .op(n27042) );
  nand2_1 U31056 ( .ip1(n27438), .ip2(\LUT[5][13] ), .op(n27041) );
  nand4_1 U31057 ( .ip1(n27044), .ip2(n27043), .ip3(n27042), .ip4(n27041), 
        .op(n27045) );
  not_ab_or_c_or_d U31058 ( .ip1(n27436), .ip2(\LUT[0][13] ), .ip3(n27046), 
        .ip4(n27045), .op(n27047) );
  nor2_1 U31059 ( .ip1(n27047), .ip2(n27446), .op(n27053) );
  nand2_1 U31060 ( .ip1(n27448), .ip2(\LUT[18][13] ), .op(n27051) );
  nand2_1 U31061 ( .ip1(n27450), .ip2(\LUT[21][13] ), .op(n27050) );
  nand2_1 U31062 ( .ip1(n27449), .ip2(\LUT[20][13] ), .op(n27049) );
  nand2_1 U31063 ( .ip1(n27451), .ip2(\LUT[16][13] ), .op(n27048) );
  nand4_1 U31064 ( .ip1(n27051), .ip2(n27050), .ip3(n27049), .ip4(n27048), 
        .op(n27052) );
  not_ab_or_c_or_d U31065 ( .ip1(\LUT[15][13] ), .ip2(n27458), .ip3(n27053), 
        .ip4(n27052), .op(n27056) );
  nand2_1 U31066 ( .ip1(n27459), .ip2(\LUT[17][13] ), .op(n27055) );
  nand2_1 U31067 ( .ip1(n27460), .ip2(\LUT[19][13] ), .op(n27054) );
  nand4_1 U31068 ( .ip1(n27057), .ip2(n27056), .ip3(n27055), .ip4(n27054), 
        .op(n27095) );
  nand2_1 U31069 ( .ip1(n27498), .ip2(\LUT[48][13] ), .op(n27061) );
  nand2_1 U31070 ( .ip1(n27499), .ip2(\LUT[49][13] ), .op(n27060) );
  nand2_1 U31071 ( .ip1(n27500), .ip2(\LUT[53][13] ), .op(n27059) );
  nand2_1 U31072 ( .ip1(n27501), .ip2(\LUT[52][13] ), .op(n27058) );
  nand4_1 U31073 ( .ip1(n27061), .ip2(n27060), .ip3(n27059), .ip4(n27058), 
        .op(n27073) );
  and2_1 U31074 ( .ip1(n27518), .ip2(\LUT[44][13] ), .op(n27067) );
  nand2_1 U31075 ( .ip1(n27507), .ip2(\LUT[54][13] ), .op(n27065) );
  nand2_1 U31076 ( .ip1(n27509), .ip2(\LUT[56][13] ), .op(n27064) );
  nand2_1 U31077 ( .ip1(n27508), .ip2(\LUT[55][13] ), .op(n27063) );
  nand2_1 U31078 ( .ip1(n27510), .ip2(\LUT[51][13] ), .op(n27062) );
  nand4_1 U31079 ( .ip1(n27065), .ip2(n27064), .ip3(n27063), .ip4(n27062), 
        .op(n27066) );
  not_ab_or_c_or_d U31080 ( .ip1(n27520), .ip2(\LUT[47][13] ), .ip3(n27067), 
        .ip4(n27066), .op(n27071) );
  nand2_1 U31081 ( .ip1(n27506), .ip2(\LUT[45][13] ), .op(n27070) );
  nand2_1 U31082 ( .ip1(n27519), .ip2(\LUT[43][13] ), .op(n27069) );
  nand2_1 U31083 ( .ip1(n27517), .ip2(\LUT[50][13] ), .op(n27068) );
  nand4_1 U31084 ( .ip1(n27071), .ip2(n27070), .ip3(n27069), .ip4(n27068), 
        .op(n27072) );
  not_ab_or_c_or_d U31085 ( .ip1(n27527), .ip2(\LUT[46][13] ), .ip3(n27073), 
        .ip4(n27072), .op(n27074) );
  nor2_1 U31086 ( .ip1(n27074), .ip2(n27528), .op(n27094) );
  nand2_1 U31087 ( .ip1(\LUT[31][13] ), .ip2(n27465), .op(n27076) );
  nand2_1 U31088 ( .ip1(\LUT[30][13] ), .ip2(n27466), .op(n27075) );
  nand2_1 U31089 ( .ip1(n27076), .ip2(n27075), .op(n27091) );
  nand2_1 U31090 ( .ip1(n27470), .ip2(\LUT[38][13] ), .op(n27080) );
  nand2_1 U31091 ( .ip1(n27469), .ip2(\LUT[39][13] ), .op(n27079) );
  nand2_1 U31092 ( .ip1(n27472), .ip2(\LUT[42][13] ), .op(n27078) );
  nand2_1 U31093 ( .ip1(n27471), .ip2(\LUT[41][13] ), .op(n27077) );
  nand4_1 U31094 ( .ip1(n27080), .ip2(n27079), .ip3(n27078), .ip4(n27077), 
        .op(n27085) );
  nand2_1 U31095 ( .ip1(\LUT[36][13] ), .ip2(n27477), .op(n27083) );
  nand2_1 U31096 ( .ip1(n27478), .ip2(\LUT[37][13] ), .op(n27082) );
  nand2_1 U31097 ( .ip1(n27479), .ip2(\LUT[32][13] ), .op(n27081) );
  nand3_1 U31098 ( .ip1(n27083), .ip2(n27082), .ip3(n27081), .op(n27084) );
  not_ab_or_c_or_d U31099 ( .ip1(n27485), .ip2(\LUT[40][13] ), .ip3(n27085), 
        .ip4(n27084), .op(n27089) );
  nand2_1 U31100 ( .ip1(n27487), .ip2(\LUT[35][13] ), .op(n27088) );
  nand2_1 U31101 ( .ip1(n27488), .ip2(\LUT[33][13] ), .op(n27087) );
  nand2_1 U31102 ( .ip1(n27486), .ip2(\LUT[34][13] ), .op(n27086) );
  nand4_1 U31103 ( .ip1(n27089), .ip2(n27088), .ip3(n27087), .ip4(n27086), 
        .op(n27090) );
  not_ab_or_c_or_d U31104 ( .ip1(n27495), .ip2(\LUT[29][13] ), .ip3(n27091), 
        .ip4(n27090), .op(n27092) );
  nor2_1 U31105 ( .ip1(n27092), .ip2(n27496), .op(n27093) );
  not_ab_or_c_or_d U31106 ( .ip1(n27533), .ip2(n27095), .ip3(n27094), .ip4(
        n27093), .op(n27096) );
  or2_1 U31107 ( .ip1(n27096), .ip2(n27265), .op(n27097) );
  nand2_1 U31108 ( .ip1(n27098), .ip2(n27097), .op(n27112) );
  nand2_1 U31109 ( .ip1(n27391), .ip2(\LUT[75][13] ), .op(n27110) );
  nand2_1 U31110 ( .ip1(n27373), .ip2(\LUT[82][13] ), .op(n27102) );
  nand2_1 U31111 ( .ip1(n27374), .ip2(\LUT[81][13] ), .op(n27101) );
  nand2_1 U31112 ( .ip1(n27375), .ip2(\LUT[84][13] ), .op(n27100) );
  nand2_1 U31113 ( .ip1(n27376), .ip2(\LUT[83][13] ), .op(n27099) );
  nand4_1 U31114 ( .ip1(n27102), .ip2(n27101), .ip3(n27100), .ip4(n27099), 
        .op(n27107) );
  nand2_1 U31115 ( .ip1(\LUT[78][13] ), .ip2(n27381), .op(n27105) );
  nand2_1 U31116 ( .ip1(n27382), .ip2(\LUT[79][13] ), .op(n27104) );
  nand2_1 U31117 ( .ip1(n27383), .ip2(\LUT[77][13] ), .op(n27103) );
  nand3_1 U31118 ( .ip1(n27105), .ip2(n27104), .ip3(n27103), .op(n27106) );
  not_ab_or_c_or_d U31119 ( .ip1(n27389), .ip2(\LUT[80][13] ), .ip3(n27107), 
        .ip4(n27106), .op(n27109) );
  nand2_1 U31120 ( .ip1(n27392), .ip2(\LUT[74][13] ), .op(n27108) );
  nand3_1 U31121 ( .ip1(n27110), .ip2(n27109), .ip3(n27108), .op(n27111) );
  not_ab_or_c_or_d U31122 ( .ip1(n27390), .ip2(\LUT[76][13] ), .ip3(n27112), 
        .ip4(n27111), .op(n27116) );
  nand2_1 U31123 ( .ip1(n27576), .ip2(\LUT[71][13] ), .op(n27115) );
  nand2_1 U31124 ( .ip1(n27569), .ip2(\LUT[73][13] ), .op(n27114) );
  nand2_1 U31125 ( .ip1(n27570), .ip2(\LUT[72][13] ), .op(n27113) );
  nand4_1 U31126 ( .ip1(n27116), .ip2(n27115), .ip3(n27114), .ip4(n27113), 
        .op(n27117) );
  nand2_1 U31127 ( .ip1(n27288), .ip2(n27117), .op(n27120) );
  nand2_1 U31128 ( .ip1(n27289), .ip2(\LUT[112][13] ), .op(n27119) );
  nand2_1 U31129 ( .ip1(n27172), .ip2(\LUT[111][13] ), .op(n27118) );
  nand4_1 U31130 ( .ip1(n27121), .ip2(n27120), .ip3(n27119), .ip4(n27118), 
        .op(n27122) );
  nand2_1 U31131 ( .ip1(n27589), .ip2(n27122), .op(n27124) );
  nand2_1 U31132 ( .ip1(sig_out[13]), .ip2(n27590), .op(n27123) );
  nand2_1 U31133 ( .ip1(n27124), .ip2(n27123), .op(n13452) );
  nand2_1 U31134 ( .ip1(n27333), .ip2(\LUT[95][14] ), .op(n27128) );
  nand2_1 U31135 ( .ip1(n27334), .ip2(\LUT[94][14] ), .op(n27127) );
  nand2_1 U31136 ( .ip1(n27335), .ip2(\LUT[98][14] ), .op(n27126) );
  nand2_1 U31137 ( .ip1(n27336), .ip2(\LUT[97][14] ), .op(n27125) );
  nand4_1 U31138 ( .ip1(n27128), .ip2(n27127), .ip3(n27126), .ip4(n27125), 
        .op(n27133) );
  nand2_1 U31139 ( .ip1(n27341), .ip2(\LUT[93][14] ), .op(n27131) );
  nand2_1 U31140 ( .ip1(n27342), .ip2(\LUT[92][14] ), .op(n27130) );
  nand2_1 U31141 ( .ip1(n27343), .ip2(\LUT[91][14] ), .op(n27129) );
  nand3_1 U31142 ( .ip1(n27131), .ip2(n27130), .ip3(n27129), .op(n27132) );
  not_ab_or_c_or_d U31143 ( .ip1(n27349), .ip2(\LUT[96][14] ), .ip3(n27133), 
        .ip4(n27132), .op(n27137) );
  nand2_1 U31144 ( .ip1(n27350), .ip2(\LUT[89][14] ), .op(n27136) );
  nand2_1 U31145 ( .ip1(n27351), .ip2(\LUT[90][14] ), .op(n27135) );
  nand2_1 U31146 ( .ip1(n27352), .ip2(\LUT[88][14] ), .op(n27134) );
  nand4_1 U31147 ( .ip1(n27137), .ip2(n27136), .ip3(n27135), .ip4(n27134), 
        .op(n27141) );
  nand2_1 U31148 ( .ip1(\LUT[85][14] ), .ip2(n27357), .op(n27139) );
  nand2_1 U31149 ( .ip1(\LUT[86][14] ), .ip2(n27358), .op(n27138) );
  nand2_1 U31150 ( .ip1(n27139), .ip2(n27138), .op(n27140) );
  not_ab_or_c_or_d U31151 ( .ip1(n27363), .ip2(\LUT[87][14] ), .ip3(n27141), 
        .ip4(n27140), .op(n27143) );
  nor2_1 U31152 ( .ip1(n27143), .ip2(n27142), .op(n27155) );
  and2_1 U31153 ( .ip1(n27317), .ip2(\LUT[105][14] ), .op(n27149) );
  nand2_1 U31154 ( .ip1(n27318), .ip2(\LUT[107][14] ), .op(n27147) );
  nand2_1 U31155 ( .ip1(n27319), .ip2(\LUT[104][14] ), .op(n27146) );
  nand2_1 U31156 ( .ip1(n27325), .ip2(\LUT[110][14] ), .op(n27145) );
  nand2_1 U31157 ( .ip1(n27309), .ip2(\LUT[109][14] ), .op(n27144) );
  nand4_1 U31158 ( .ip1(n27147), .ip2(n27146), .ip3(n27145), .ip4(n27144), 
        .op(n27148) );
  not_ab_or_c_or_d U31159 ( .ip1(\LUT[102][14] ), .ip2(n27326), .ip3(n27149), 
        .ip4(n27148), .op(n27153) );
  nand2_1 U31160 ( .ip1(n27370), .ip2(\LUT[100][14] ), .op(n27152) );
  nand2_1 U31161 ( .ip1(n27328), .ip2(\LUT[101][14] ), .op(n27151) );
  nand2_1 U31162 ( .ip1(n27327), .ip2(\LUT[103][14] ), .op(n27150) );
  nand4_1 U31163 ( .ip1(n27153), .ip2(n27152), .ip3(n27151), .ip4(n27150), 
        .op(n27154) );
  not_ab_or_c_or_d U31164 ( .ip1(\LUT[99][14] ), .ip2(n27156), .ip3(n27155), 
        .ip4(n27154), .op(n27157) );
  nor2_1 U31165 ( .ip1(n27157), .ip2(n27371), .op(n27171) );
  nand2_1 U31166 ( .ip1(n27582), .ip2(\LUT[115][14] ), .op(n27161) );
  nand2_1 U31167 ( .ip1(n27298), .ip2(\LUT[117][14] ), .op(n27160) );
  nand2_1 U31168 ( .ip1(n27299), .ip2(\LUT[118][14] ), .op(n27159) );
  nand2_1 U31169 ( .ip1(n27300), .ip2(\LUT[119][14] ), .op(n27158) );
  nand4_1 U31170 ( .ip1(n27161), .ip2(n27160), .ip3(n27159), .ip4(n27158), 
        .op(n27162) );
  or2_1 U31171 ( .ip1(n27297), .ip2(n27162), .op(n27164) );
  or2_1 U31172 ( .ip1(\LUT[116][14] ), .ip2(n27162), .op(n27163) );
  nand2_1 U31173 ( .ip1(n27164), .ip2(n27163), .op(n27169) );
  nand2_1 U31174 ( .ip1(n27583), .ip2(\LUT[113][14] ), .op(n27168) );
  nand2_1 U31175 ( .ip1(n27165), .ip2(\LUT[108][14] ), .op(n27167) );
  nand2_1 U31176 ( .ip1(n27305), .ip2(\LUT[114][14] ), .op(n27166) );
  nand4_1 U31177 ( .ip1(n27169), .ip2(n27168), .ip3(n27167), .ip4(n27166), 
        .op(n27170) );
  not_ab_or_c_or_d U31178 ( .ip1(n27172), .ip2(\LUT[111][14] ), .ip3(n27171), 
        .ip4(n27170), .op(n27293) );
  and2_1 U31179 ( .ip1(n27548), .ip2(\LUT[67][14] ), .op(n27178) );
  nand2_1 U31180 ( .ip1(n27534), .ip2(\LUT[65][14] ), .op(n27176) );
  nand2_1 U31181 ( .ip1(n27537), .ip2(\LUT[68][14] ), .op(n27175) );
  nand2_1 U31182 ( .ip1(n27535), .ip2(\LUT[69][14] ), .op(n27174) );
  nand2_1 U31183 ( .ip1(n27536), .ip2(\LUT[70][14] ), .op(n27173) );
  nand4_1 U31184 ( .ip1(n27176), .ip2(n27175), .ip3(n27174), .ip4(n27173), 
        .op(n27177) );
  not_ab_or_c_or_d U31185 ( .ip1(n27542), .ip2(\LUT[66][14] ), .ip3(n27178), 
        .ip4(n27177), .op(n27182) );
  nand2_1 U31186 ( .ip1(n27546), .ip2(\LUT[59][14] ), .op(n27181) );
  nand2_1 U31187 ( .ip1(n27556), .ip2(\LUT[63][14] ), .op(n27180) );
  nand2_1 U31188 ( .ip1(n27547), .ip2(\LUT[64][14] ), .op(n27179) );
  nand4_1 U31189 ( .ip1(n27182), .ip2(n27181), .ip3(n27180), .ip4(n27179), 
        .op(n27188) );
  nand2_1 U31190 ( .ip1(n27397), .ip2(\LUT[58][14] ), .op(n27186) );
  nand2_1 U31191 ( .ip1(n27554), .ip2(\LUT[60][14] ), .op(n27185) );
  nand2_1 U31192 ( .ip1(n27555), .ip2(\LUT[61][14] ), .op(n27184) );
  nand2_1 U31193 ( .ip1(n27563), .ip2(\LUT[62][14] ), .op(n27183) );
  nand4_1 U31194 ( .ip1(n27186), .ip2(n27185), .ip3(n27184), .ip4(n27183), 
        .op(n27187) );
  not_ab_or_c_or_d U31195 ( .ip1(n27553), .ip2(\LUT[57][14] ), .ip3(n27188), 
        .ip4(n27187), .op(n27189) );
  or2_1 U31196 ( .ip1(n27189), .ip2(n27265), .op(n27268) );
  nand2_1 U31197 ( .ip1(\LUT[27][14] ), .ip2(n27398), .op(n27192) );
  nand2_1 U31198 ( .ip1(n27399), .ip2(\LUT[26][14] ), .op(n27191) );
  nand2_1 U31199 ( .ip1(n27400), .ip2(\LUT[28][14] ), .op(n27190) );
  nand3_1 U31200 ( .ip1(n27192), .ip2(n27191), .ip3(n27190), .op(n27197) );
  nand2_1 U31201 ( .ip1(\LUT[24][14] ), .ip2(n27404), .op(n27195) );
  nand2_1 U31202 ( .ip1(n27405), .ip2(\LUT[25][14] ), .op(n27194) );
  nand2_1 U31203 ( .ip1(n27406), .ip2(\LUT[23][14] ), .op(n27193) );
  nand3_1 U31204 ( .ip1(n27195), .ip2(n27194), .ip3(n27193), .op(n27196) );
  not_ab_or_c_or_d U31205 ( .ip1(n27460), .ip2(\LUT[19][14] ), .ip3(n27197), 
        .ip4(n27196), .op(n27226) );
  nand2_1 U31206 ( .ip1(\LUT[2][14] ), .ip2(n27413), .op(n27199) );
  nand2_1 U31207 ( .ip1(\LUT[3][14] ), .ip2(n27414), .op(n27198) );
  nand2_1 U31208 ( .ip1(n27199), .ip2(n27198), .op(n27215) );
  nand2_1 U31209 ( .ip1(n27417), .ip2(\LUT[7][14] ), .op(n27203) );
  nand2_1 U31210 ( .ip1(n27427), .ip2(\LUT[12][14] ), .op(n27202) );
  nand2_1 U31211 ( .ip1(n27419), .ip2(\LUT[14][14] ), .op(n27201) );
  nand2_1 U31212 ( .ip1(n27420), .ip2(\LUT[13][14] ), .op(n27200) );
  nand4_1 U31213 ( .ip1(n27203), .ip2(n27202), .ip3(n27201), .ip4(n27200), 
        .op(n27209) );
  nand2_1 U31214 ( .ip1(n27426), .ip2(\LUT[8][14] ), .op(n27207) );
  nand2_1 U31215 ( .ip1(n27435), .ip2(\LUT[11][14] ), .op(n27206) );
  nand2_1 U31216 ( .ip1(n27425), .ip2(\LUT[10][14] ), .op(n27205) );
  nand2_1 U31217 ( .ip1(n27428), .ip2(\LUT[6][14] ), .op(n27204) );
  nand4_1 U31218 ( .ip1(n27207), .ip2(n27206), .ip3(n27205), .ip4(n27204), 
        .op(n27208) );
  not_ab_or_c_or_d U31219 ( .ip1(n27418), .ip2(\LUT[9][14] ), .ip3(n27209), 
        .ip4(n27208), .op(n27213) );
  nand2_1 U31220 ( .ip1(n27436), .ip2(\LUT[0][14] ), .op(n27212) );
  nand2_1 U31221 ( .ip1(n27438), .ip2(\LUT[5][14] ), .op(n27211) );
  nand2_1 U31222 ( .ip1(n27437), .ip2(\LUT[4][14] ), .op(n27210) );
  nand4_1 U31223 ( .ip1(n27213), .ip2(n27212), .ip3(n27211), .ip4(n27210), 
        .op(n27214) );
  not_ab_or_c_or_d U31224 ( .ip1(n27445), .ip2(\LUT[1][14] ), .ip3(n27215), 
        .ip4(n27214), .op(n27216) );
  nor2_1 U31225 ( .ip1(n27216), .ip2(n27446), .op(n27222) );
  nand2_1 U31226 ( .ip1(n27450), .ip2(\LUT[21][14] ), .op(n27220) );
  nand2_1 U31227 ( .ip1(n27449), .ip2(\LUT[20][14] ), .op(n27219) );
  nand2_1 U31228 ( .ip1(n27448), .ip2(\LUT[18][14] ), .op(n27218) );
  nand2_1 U31229 ( .ip1(n27451), .ip2(\LUT[16][14] ), .op(n27217) );
  nand4_1 U31230 ( .ip1(n27220), .ip2(n27219), .ip3(n27218), .ip4(n27217), 
        .op(n27221) );
  not_ab_or_c_or_d U31231 ( .ip1(\LUT[15][14] ), .ip2(n27458), .ip3(n27222), 
        .ip4(n27221), .op(n27225) );
  nand2_1 U31232 ( .ip1(n27412), .ip2(\LUT[22][14] ), .op(n27224) );
  nand2_1 U31233 ( .ip1(n27459), .ip2(\LUT[17][14] ), .op(n27223) );
  nand4_1 U31234 ( .ip1(n27226), .ip2(n27225), .ip3(n27224), .ip4(n27223), 
        .op(n27264) );
  nand2_1 U31235 ( .ip1(\LUT[31][14] ), .ip2(n27465), .op(n27228) );
  nand2_1 U31236 ( .ip1(\LUT[30][14] ), .ip2(n27466), .op(n27227) );
  nand2_1 U31237 ( .ip1(n27228), .ip2(n27227), .op(n27243) );
  nand2_1 U31238 ( .ip1(n27470), .ip2(\LUT[38][14] ), .op(n27232) );
  nand2_1 U31239 ( .ip1(n27469), .ip2(\LUT[39][14] ), .op(n27231) );
  nand2_1 U31240 ( .ip1(n27472), .ip2(\LUT[42][14] ), .op(n27230) );
  nand2_1 U31241 ( .ip1(n27471), .ip2(\LUT[41][14] ), .op(n27229) );
  nand4_1 U31242 ( .ip1(n27232), .ip2(n27231), .ip3(n27230), .ip4(n27229), 
        .op(n27237) );
  nand2_1 U31243 ( .ip1(\LUT[36][14] ), .ip2(n27477), .op(n27235) );
  nand2_1 U31244 ( .ip1(n27478), .ip2(\LUT[37][14] ), .op(n27234) );
  nand2_1 U31245 ( .ip1(n27488), .ip2(\LUT[33][14] ), .op(n27233) );
  nand3_1 U31246 ( .ip1(n27235), .ip2(n27234), .ip3(n27233), .op(n27236) );
  not_ab_or_c_or_d U31247 ( .ip1(n27485), .ip2(\LUT[40][14] ), .ip3(n27237), 
        .ip4(n27236), .op(n27241) );
  nand2_1 U31248 ( .ip1(n27479), .ip2(\LUT[32][14] ), .op(n27240) );
  nand2_1 U31249 ( .ip1(n27486), .ip2(\LUT[34][14] ), .op(n27239) );
  nand2_1 U31250 ( .ip1(n27487), .ip2(\LUT[35][14] ), .op(n27238) );
  nand4_1 U31251 ( .ip1(n27241), .ip2(n27240), .ip3(n27239), .ip4(n27238), 
        .op(n27242) );
  not_ab_or_c_or_d U31252 ( .ip1(n27495), .ip2(\LUT[29][14] ), .ip3(n27243), 
        .ip4(n27242), .op(n27244) );
  nor2_1 U31253 ( .ip1(n27244), .ip2(n27496), .op(n27263) );
  nand2_1 U31254 ( .ip1(n27498), .ip2(\LUT[48][14] ), .op(n27248) );
  nand2_1 U31255 ( .ip1(n27499), .ip2(\LUT[49][14] ), .op(n27247) );
  nand2_1 U31256 ( .ip1(n27507), .ip2(\LUT[54][14] ), .op(n27246) );
  nand2_1 U31257 ( .ip1(n27501), .ip2(\LUT[52][14] ), .op(n27245) );
  nand4_1 U31258 ( .ip1(n27248), .ip2(n27247), .ip3(n27246), .ip4(n27245), 
        .op(n27260) );
  and2_1 U31259 ( .ip1(n27506), .ip2(\LUT[45][14] ), .op(n27254) );
  nand2_1 U31260 ( .ip1(n27509), .ip2(\LUT[56][14] ), .op(n27252) );
  nand2_1 U31261 ( .ip1(n27510), .ip2(\LUT[51][14] ), .op(n27251) );
  nand2_1 U31262 ( .ip1(n27508), .ip2(\LUT[55][14] ), .op(n27250) );
  nand2_1 U31263 ( .ip1(n27500), .ip2(\LUT[53][14] ), .op(n27249) );
  nand4_1 U31264 ( .ip1(n27252), .ip2(n27251), .ip3(n27250), .ip4(n27249), 
        .op(n27253) );
  not_ab_or_c_or_d U31265 ( .ip1(n27517), .ip2(\LUT[50][14] ), .ip3(n27254), 
        .ip4(n27253), .op(n27258) );
  nand2_1 U31266 ( .ip1(n27518), .ip2(\LUT[44][14] ), .op(n27257) );
  nand2_1 U31267 ( .ip1(n27519), .ip2(\LUT[43][14] ), .op(n27256) );
  nand2_1 U31268 ( .ip1(n27520), .ip2(\LUT[47][14] ), .op(n27255) );
  nand4_1 U31269 ( .ip1(n27258), .ip2(n27257), .ip3(n27256), .ip4(n27255), 
        .op(n27259) );
  not_ab_or_c_or_d U31270 ( .ip1(n27527), .ip2(\LUT[46][14] ), .ip3(n27260), 
        .ip4(n27259), .op(n27261) );
  nor2_1 U31271 ( .ip1(n27261), .ip2(n27528), .op(n27262) );
  not_ab_or_c_or_d U31272 ( .ip1(n27533), .ip2(n27264), .ip3(n27263), .ip4(
        n27262), .op(n27266) );
  or2_1 U31273 ( .ip1(n27266), .ip2(n27265), .op(n27267) );
  nand2_1 U31274 ( .ip1(n27268), .ip2(n27267), .op(n27282) );
  nand2_1 U31275 ( .ip1(n27391), .ip2(\LUT[75][14] ), .op(n27280) );
  nand2_1 U31276 ( .ip1(n27373), .ip2(\LUT[82][14] ), .op(n27272) );
  nand2_1 U31277 ( .ip1(n27374), .ip2(\LUT[81][14] ), .op(n27271) );
  nand2_1 U31278 ( .ip1(n27375), .ip2(\LUT[84][14] ), .op(n27270) );
  nand2_1 U31279 ( .ip1(n27376), .ip2(\LUT[83][14] ), .op(n27269) );
  nand4_1 U31280 ( .ip1(n27272), .ip2(n27271), .ip3(n27270), .ip4(n27269), 
        .op(n27277) );
  nand2_1 U31281 ( .ip1(\LUT[78][14] ), .ip2(n27381), .op(n27275) );
  nand2_1 U31282 ( .ip1(n27382), .ip2(\LUT[79][14] ), .op(n27274) );
  nand2_1 U31283 ( .ip1(n27383), .ip2(\LUT[77][14] ), .op(n27273) );
  nand3_1 U31284 ( .ip1(n27275), .ip2(n27274), .ip3(n27273), .op(n27276) );
  not_ab_or_c_or_d U31285 ( .ip1(n27389), .ip2(\LUT[80][14] ), .ip3(n27277), 
        .ip4(n27276), .op(n27279) );
  nand2_1 U31286 ( .ip1(n27392), .ip2(\LUT[74][14] ), .op(n27278) );
  nand3_1 U31287 ( .ip1(n27280), .ip2(n27279), .ip3(n27278), .op(n27281) );
  not_ab_or_c_or_d U31288 ( .ip1(n27390), .ip2(\LUT[76][14] ), .ip3(n27282), 
        .ip4(n27281), .op(n27286) );
  nand2_1 U31289 ( .ip1(n27576), .ip2(\LUT[71][14] ), .op(n27285) );
  nand2_1 U31290 ( .ip1(n27570), .ip2(\LUT[72][14] ), .op(n27284) );
  nand2_1 U31291 ( .ip1(n27569), .ip2(\LUT[73][14] ), .op(n27283) );
  nand4_1 U31292 ( .ip1(n27286), .ip2(n27285), .ip3(n27284), .ip4(n27283), 
        .op(n27287) );
  nand2_1 U31293 ( .ip1(n27288), .ip2(n27287), .op(n27292) );
  nand2_1 U31294 ( .ip1(n27581), .ip2(\LUT[106][14] ), .op(n27291) );
  nand2_1 U31295 ( .ip1(n27289), .ip2(\LUT[112][14] ), .op(n27290) );
  nand4_1 U31296 ( .ip1(n27293), .ip2(n27292), .ip3(n27291), .ip4(n27290), 
        .op(n27294) );
  nand2_1 U31297 ( .ip1(n27589), .ip2(n27294), .op(n27296) );
  nand2_1 U31298 ( .ip1(sig_out[14]), .ip2(n27590), .op(n27295) );
  nand2_1 U31299 ( .ip1(n27296), .ip2(n27295), .op(n13451) );
  nand2_1 U31300 ( .ip1(n27297), .ip2(\LUT[116][15] ), .op(n27304) );
  nand2_1 U31301 ( .ip1(n27298), .ip2(\LUT[117][15] ), .op(n27303) );
  nand2_1 U31302 ( .ip1(n27299), .ip2(\LUT[118][15] ), .op(n27302) );
  nand2_1 U31303 ( .ip1(n27300), .ip2(\LUT[119][15] ), .op(n27301) );
  nand4_1 U31304 ( .ip1(n27304), .ip2(n27303), .ip3(n27302), .ip4(n27301), 
        .op(n27306) );
  or2_1 U31305 ( .ip1(n27305), .ip2(n27306), .op(n27308) );
  or2_1 U31306 ( .ip1(\LUT[114][15] ), .ip2(n27306), .op(n27307) );
  nand2_1 U31307 ( .ip1(n27308), .ip2(n27307), .op(n27587) );
  nand2_1 U31308 ( .ip1(n27309), .ip2(\LUT[109][15] ), .op(n27316) );
  nand2_1 U31309 ( .ip1(n27310), .ip2(\LUT[108][15] ), .op(n27315) );
  nand2_1 U31310 ( .ip1(n27311), .ip2(\LUT[111][15] ), .op(n27314) );
  nand2_1 U31311 ( .ip1(n27312), .ip2(\LUT[112][15] ), .op(n27313) );
  nand4_1 U31312 ( .ip1(n27316), .ip2(n27315), .ip3(n27314), .ip4(n27313), 
        .op(n27324) );
  nand2_1 U31313 ( .ip1(\LUT[105][15] ), .ip2(n27317), .op(n27322) );
  nand2_1 U31314 ( .ip1(n27318), .ip2(\LUT[107][15] ), .op(n27321) );
  nand2_1 U31315 ( .ip1(n27319), .ip2(\LUT[104][15] ), .op(n27320) );
  nand3_1 U31316 ( .ip1(n27322), .ip2(n27321), .ip3(n27320), .op(n27323) );
  not_ab_or_c_or_d U31317 ( .ip1(n27325), .ip2(\LUT[110][15] ), .ip3(n27324), 
        .ip4(n27323), .op(n27332) );
  nand2_1 U31318 ( .ip1(n27326), .ip2(\LUT[102][15] ), .op(n27331) );
  nand2_1 U31319 ( .ip1(n27327), .ip2(\LUT[103][15] ), .op(n27330) );
  nand2_1 U31320 ( .ip1(n27328), .ip2(\LUT[101][15] ), .op(n27329) );
  nand4_1 U31321 ( .ip1(n27332), .ip2(n27331), .ip3(n27330), .ip4(n27329), 
        .op(n27369) );
  nand2_1 U31322 ( .ip1(n27333), .ip2(\LUT[95][15] ), .op(n27340) );
  nand2_1 U31323 ( .ip1(n27334), .ip2(\LUT[94][15] ), .op(n27339) );
  nand2_1 U31324 ( .ip1(n27335), .ip2(\LUT[98][15] ), .op(n27338) );
  nand2_1 U31325 ( .ip1(n27336), .ip2(\LUT[97][15] ), .op(n27337) );
  nand4_1 U31326 ( .ip1(n27340), .ip2(n27339), .ip3(n27338), .ip4(n27337), 
        .op(n27348) );
  nand2_1 U31327 ( .ip1(n27341), .ip2(\LUT[93][15] ), .op(n27346) );
  nand2_1 U31328 ( .ip1(n27342), .ip2(\LUT[92][15] ), .op(n27345) );
  nand2_1 U31329 ( .ip1(n27343), .ip2(\LUT[91][15] ), .op(n27344) );
  nand3_1 U31330 ( .ip1(n27346), .ip2(n27345), .ip3(n27344), .op(n27347) );
  not_ab_or_c_or_d U31331 ( .ip1(n27349), .ip2(\LUT[96][15] ), .ip3(n27348), 
        .ip4(n27347), .op(n27356) );
  nand2_1 U31332 ( .ip1(n27350), .ip2(\LUT[89][15] ), .op(n27355) );
  nand2_1 U31333 ( .ip1(n27351), .ip2(\LUT[90][15] ), .op(n27354) );
  nand2_1 U31334 ( .ip1(n27352), .ip2(\LUT[88][15] ), .op(n27353) );
  nand4_1 U31335 ( .ip1(n27356), .ip2(n27355), .ip3(n27354), .ip4(n27353), 
        .op(n27362) );
  nand2_1 U31336 ( .ip1(\LUT[85][15] ), .ip2(n27357), .op(n27360) );
  nand2_1 U31337 ( .ip1(\LUT[86][15] ), .ip2(n27358), .op(n27359) );
  nand2_1 U31338 ( .ip1(n27360), .ip2(n27359), .op(n27361) );
  not_ab_or_c_or_d U31339 ( .ip1(n27363), .ip2(\LUT[87][15] ), .ip3(n27362), 
        .ip4(n27361), .op(n27366) );
  nor2_1 U31340 ( .ip1(\LUT[99][15] ), .ip2(n27367), .op(n27365) );
  not_ab_or_c_or_d U31341 ( .ip1(n27367), .ip2(n27366), .ip3(n27365), .ip4(
        n27364), .op(n27368) );
  not_ab_or_c_or_d U31342 ( .ip1(n27370), .ip2(\LUT[100][15] ), .ip3(n27369), 
        .ip4(n27368), .op(n27372) );
  nor2_1 U31343 ( .ip1(n27372), .ip2(n27371), .op(n27580) );
  nand2_1 U31344 ( .ip1(n27373), .ip2(\LUT[82][15] ), .op(n27380) );
  nand2_1 U31345 ( .ip1(n27374), .ip2(\LUT[81][15] ), .op(n27379) );
  nand2_1 U31346 ( .ip1(n27375), .ip2(\LUT[84][15] ), .op(n27378) );
  nand2_1 U31347 ( .ip1(n27376), .ip2(\LUT[83][15] ), .op(n27377) );
  nand4_1 U31348 ( .ip1(n27380), .ip2(n27379), .ip3(n27378), .ip4(n27377), 
        .op(n27388) );
  nand2_1 U31349 ( .ip1(\LUT[78][15] ), .ip2(n27381), .op(n27386) );
  nand2_1 U31350 ( .ip1(n27382), .ip2(\LUT[79][15] ), .op(n27385) );
  nand2_1 U31351 ( .ip1(n27383), .ip2(\LUT[77][15] ), .op(n27384) );
  nand3_1 U31352 ( .ip1(n27386), .ip2(n27385), .ip3(n27384), .op(n27387) );
  not_ab_or_c_or_d U31353 ( .ip1(n27389), .ip2(\LUT[80][15] ), .ip3(n27388), 
        .ip4(n27387), .op(n27396) );
  nand2_1 U31354 ( .ip1(n27390), .ip2(\LUT[76][15] ), .op(n27395) );
  nand2_1 U31355 ( .ip1(n27391), .ip2(\LUT[75][15] ), .op(n27394) );
  nand2_1 U31356 ( .ip1(n27392), .ip2(\LUT[74][15] ), .op(n27393) );
  nand4_1 U31357 ( .ip1(n27396), .ip2(n27395), .ip3(n27394), .ip4(n27393), 
        .op(n27575) );
  nand2_1 U31358 ( .ip1(\LUT[58][15] ), .ip2(n27397), .op(n27566) );
  nand2_1 U31359 ( .ip1(\LUT[27][15] ), .ip2(n27398), .op(n27403) );
  nand2_1 U31360 ( .ip1(n27399), .ip2(\LUT[26][15] ), .op(n27402) );
  nand2_1 U31361 ( .ip1(n27400), .ip2(\LUT[28][15] ), .op(n27401) );
  nand3_1 U31362 ( .ip1(n27403), .ip2(n27402), .ip3(n27401), .op(n27411) );
  nand2_1 U31363 ( .ip1(n27404), .ip2(\LUT[24][15] ), .op(n27409) );
  nand2_1 U31364 ( .ip1(n27405), .ip2(\LUT[25][15] ), .op(n27408) );
  nand2_1 U31365 ( .ip1(n27406), .ip2(\LUT[23][15] ), .op(n27407) );
  nand3_1 U31366 ( .ip1(n27409), .ip2(n27408), .ip3(n27407), .op(n27410) );
  not_ab_or_c_or_d U31367 ( .ip1(n27412), .ip2(\LUT[22][15] ), .ip3(n27411), 
        .ip4(n27410), .op(n27464) );
  nand2_1 U31368 ( .ip1(\LUT[2][15] ), .ip2(n27413), .op(n27416) );
  nand2_1 U31369 ( .ip1(\LUT[3][15] ), .ip2(n27414), .op(n27415) );
  nand2_1 U31370 ( .ip1(n27416), .ip2(n27415), .op(n27444) );
  nand2_1 U31371 ( .ip1(n27417), .ip2(\LUT[7][15] ), .op(n27424) );
  nand2_1 U31372 ( .ip1(n27418), .ip2(\LUT[9][15] ), .op(n27423) );
  nand2_1 U31373 ( .ip1(n27419), .ip2(\LUT[14][15] ), .op(n27422) );
  nand2_1 U31374 ( .ip1(n27420), .ip2(\LUT[13][15] ), .op(n27421) );
  nand4_1 U31375 ( .ip1(n27424), .ip2(n27423), .ip3(n27422), .ip4(n27421), 
        .op(n27434) );
  nand2_1 U31376 ( .ip1(n27425), .ip2(\LUT[10][15] ), .op(n27432) );
  nand2_1 U31377 ( .ip1(n27426), .ip2(\LUT[8][15] ), .op(n27431) );
  nand2_1 U31378 ( .ip1(n27427), .ip2(\LUT[12][15] ), .op(n27430) );
  nand2_1 U31379 ( .ip1(n27428), .ip2(\LUT[6][15] ), .op(n27429) );
  nand4_1 U31380 ( .ip1(n27432), .ip2(n27431), .ip3(n27430), .ip4(n27429), 
        .op(n27433) );
  not_ab_or_c_or_d U31381 ( .ip1(n27435), .ip2(\LUT[11][15] ), .ip3(n27434), 
        .ip4(n27433), .op(n27442) );
  nand2_1 U31382 ( .ip1(n27436), .ip2(\LUT[0][15] ), .op(n27441) );
  nand2_1 U31383 ( .ip1(n27437), .ip2(\LUT[4][15] ), .op(n27440) );
  nand2_1 U31384 ( .ip1(n27438), .ip2(\LUT[5][15] ), .op(n27439) );
  nand4_1 U31385 ( .ip1(n27442), .ip2(n27441), .ip3(n27440), .ip4(n27439), 
        .op(n27443) );
  not_ab_or_c_or_d U31386 ( .ip1(n27445), .ip2(\LUT[1][15] ), .ip3(n27444), 
        .ip4(n27443), .op(n27447) );
  nor2_1 U31387 ( .ip1(n27447), .ip2(n27446), .op(n27457) );
  nand2_1 U31388 ( .ip1(n27448), .ip2(\LUT[18][15] ), .op(n27455) );
  nand2_1 U31389 ( .ip1(n27449), .ip2(\LUT[20][15] ), .op(n27454) );
  nand2_1 U31390 ( .ip1(n27450), .ip2(\LUT[21][15] ), .op(n27453) );
  nand2_1 U31391 ( .ip1(n27451), .ip2(\LUT[16][15] ), .op(n27452) );
  nand4_1 U31392 ( .ip1(n27455), .ip2(n27454), .ip3(n27453), .ip4(n27452), 
        .op(n27456) );
  not_ab_or_c_or_d U31393 ( .ip1(\LUT[15][15] ), .ip2(n27458), .ip3(n27457), 
        .ip4(n27456), .op(n27463) );
  nand2_1 U31394 ( .ip1(n27459), .ip2(\LUT[17][15] ), .op(n27462) );
  nand2_1 U31395 ( .ip1(n27460), .ip2(\LUT[19][15] ), .op(n27461) );
  nand4_1 U31396 ( .ip1(n27464), .ip2(n27463), .ip3(n27462), .ip4(n27461), 
        .op(n27532) );
  nand2_1 U31397 ( .ip1(\LUT[31][15] ), .ip2(n27465), .op(n27468) );
  nand2_1 U31398 ( .ip1(\LUT[30][15] ), .ip2(n27466), .op(n27467) );
  nand2_1 U31399 ( .ip1(n27468), .ip2(n27467), .op(n27494) );
  nand2_1 U31400 ( .ip1(n27469), .ip2(\LUT[39][15] ), .op(n27476) );
  nand2_1 U31401 ( .ip1(n27470), .ip2(\LUT[38][15] ), .op(n27475) );
  nand2_1 U31402 ( .ip1(n27471), .ip2(\LUT[41][15] ), .op(n27474) );
  nand2_1 U31403 ( .ip1(n27472), .ip2(\LUT[42][15] ), .op(n27473) );
  nand4_1 U31404 ( .ip1(n27476), .ip2(n27475), .ip3(n27474), .ip4(n27473), 
        .op(n27484) );
  nand2_1 U31405 ( .ip1(\LUT[36][15] ), .ip2(n27477), .op(n27482) );
  nand2_1 U31406 ( .ip1(n27478), .ip2(\LUT[37][15] ), .op(n27481) );
  nand2_1 U31407 ( .ip1(n27479), .ip2(\LUT[32][15] ), .op(n27480) );
  nand3_1 U31408 ( .ip1(n27482), .ip2(n27481), .ip3(n27480), .op(n27483) );
  not_ab_or_c_or_d U31409 ( .ip1(n27485), .ip2(\LUT[40][15] ), .ip3(n27484), 
        .ip4(n27483), .op(n27492) );
  nand2_1 U31410 ( .ip1(n27486), .ip2(\LUT[34][15] ), .op(n27491) );
  nand2_1 U31411 ( .ip1(n27487), .ip2(\LUT[35][15] ), .op(n27490) );
  nand2_1 U31412 ( .ip1(n27488), .ip2(\LUT[33][15] ), .op(n27489) );
  nand4_1 U31413 ( .ip1(n27492), .ip2(n27491), .ip3(n27490), .ip4(n27489), 
        .op(n27493) );
  not_ab_or_c_or_d U31414 ( .ip1(n27495), .ip2(\LUT[29][15] ), .ip3(n27494), 
        .ip4(n27493), .op(n27497) );
  nor2_1 U31415 ( .ip1(n27497), .ip2(n27496), .op(n27531) );
  nand2_1 U31416 ( .ip1(n27498), .ip2(\LUT[48][15] ), .op(n27505) );
  nand2_1 U31417 ( .ip1(n27499), .ip2(\LUT[49][15] ), .op(n27504) );
  nand2_1 U31418 ( .ip1(n27500), .ip2(\LUT[53][15] ), .op(n27503) );
  nand2_1 U31419 ( .ip1(n27501), .ip2(\LUT[52][15] ), .op(n27502) );
  nand4_1 U31420 ( .ip1(n27505), .ip2(n27504), .ip3(n27503), .ip4(n27502), 
        .op(n27526) );
  and2_1 U31421 ( .ip1(n27506), .ip2(\LUT[45][15] ), .op(n27516) );
  nand2_1 U31422 ( .ip1(n27507), .ip2(\LUT[54][15] ), .op(n27514) );
  nand2_1 U31423 ( .ip1(n27508), .ip2(\LUT[55][15] ), .op(n27513) );
  nand2_1 U31424 ( .ip1(n27509), .ip2(\LUT[56][15] ), .op(n27512) );
  nand2_1 U31425 ( .ip1(n27510), .ip2(\LUT[51][15] ), .op(n27511) );
  nand4_1 U31426 ( .ip1(n27514), .ip2(n27513), .ip3(n27512), .ip4(n27511), 
        .op(n27515) );
  not_ab_or_c_or_d U31427 ( .ip1(n27517), .ip2(\LUT[50][15] ), .ip3(n27516), 
        .ip4(n27515), .op(n27524) );
  nand2_1 U31428 ( .ip1(n27518), .ip2(\LUT[44][15] ), .op(n27523) );
  nand2_1 U31429 ( .ip1(n27519), .ip2(\LUT[43][15] ), .op(n27522) );
  nand2_1 U31430 ( .ip1(n27520), .ip2(\LUT[47][15] ), .op(n27521) );
  nand4_1 U31431 ( .ip1(n27524), .ip2(n27523), .ip3(n27522), .ip4(n27521), 
        .op(n27525) );
  not_ab_or_c_or_d U31432 ( .ip1(n27527), .ip2(\LUT[46][15] ), .ip3(n27526), 
        .ip4(n27525), .op(n27529) );
  nor2_1 U31433 ( .ip1(n27529), .ip2(n27528), .op(n27530) );
  not_ab_or_c_or_d U31434 ( .ip1(n27533), .ip2(n27532), .ip3(n27531), .ip4(
        n27530), .op(n27565) );
  nand2_1 U31435 ( .ip1(n27534), .ip2(\LUT[65][15] ), .op(n27541) );
  nand2_1 U31436 ( .ip1(n27535), .ip2(\LUT[69][15] ), .op(n27540) );
  nand2_1 U31437 ( .ip1(n27536), .ip2(\LUT[70][15] ), .op(n27539) );
  nand2_1 U31438 ( .ip1(n27537), .ip2(\LUT[68][15] ), .op(n27538) );
  nand4_1 U31439 ( .ip1(n27541), .ip2(n27540), .ip3(n27539), .ip4(n27538), 
        .op(n27543) );
  or2_1 U31440 ( .ip1(n27542), .ip2(n27543), .op(n27545) );
  or2_1 U31441 ( .ip1(\LUT[66][15] ), .ip2(n27543), .op(n27544) );
  nand2_1 U31442 ( .ip1(n27545), .ip2(n27544), .op(n27552) );
  nand2_1 U31443 ( .ip1(n27546), .ip2(\LUT[59][15] ), .op(n27551) );
  nand2_1 U31444 ( .ip1(n27547), .ip2(\LUT[64][15] ), .op(n27550) );
  nand2_1 U31445 ( .ip1(n27548), .ip2(\LUT[67][15] ), .op(n27549) );
  nand4_1 U31446 ( .ip1(n27552), .ip2(n27551), .ip3(n27550), .ip4(n27549), 
        .op(n27562) );
  nand2_1 U31447 ( .ip1(n27553), .ip2(\LUT[57][15] ), .op(n27560) );
  nand2_1 U31448 ( .ip1(n27554), .ip2(\LUT[60][15] ), .op(n27559) );
  nand2_1 U31449 ( .ip1(n27555), .ip2(\LUT[61][15] ), .op(n27558) );
  nand2_1 U31450 ( .ip1(n27556), .ip2(\LUT[63][15] ), .op(n27557) );
  nand4_1 U31451 ( .ip1(n27560), .ip2(n27559), .ip3(n27558), .ip4(n27557), 
        .op(n27561) );
  not_ab_or_c_or_d U31452 ( .ip1(n27563), .ip2(\LUT[62][15] ), .ip3(n27562), 
        .ip4(n27561), .op(n27564) );
  nand3_1 U31453 ( .ip1(n27566), .ip2(n27565), .ip3(n27564), .op(n27568) );
  nand2_1 U31454 ( .ip1(n27568), .ip2(n27567), .op(n27573) );
  nand2_1 U31455 ( .ip1(n27569), .ip2(\LUT[73][15] ), .op(n27572) );
  nand2_1 U31456 ( .ip1(n27570), .ip2(\LUT[72][15] ), .op(n27571) );
  nand3_1 U31457 ( .ip1(n27573), .ip2(n27572), .ip3(n27571), .op(n27574) );
  not_ab_or_c_or_d U31458 ( .ip1(n27576), .ip2(\LUT[71][15] ), .ip3(n27575), 
        .ip4(n27574), .op(n27578) );
  nor2_1 U31459 ( .ip1(n27578), .ip2(n27577), .op(n27579) );
  not_ab_or_c_or_d U31460 ( .ip1(n27581), .ip2(\LUT[106][15] ), .ip3(n27580), 
        .ip4(n27579), .op(n27586) );
  nand2_1 U31461 ( .ip1(n27582), .ip2(\LUT[115][15] ), .op(n27585) );
  nand2_1 U31462 ( .ip1(n27583), .ip2(\LUT[113][15] ), .op(n27584) );
  nand4_1 U31463 ( .ip1(n27587), .ip2(n27586), .ip3(n27585), .ip4(n27584), 
        .op(n27588) );
  nand2_1 U31464 ( .ip1(n27589), .ip2(n27588), .op(n27592) );
  nand2_1 U31465 ( .ip1(sig_out[15]), .ip2(n27590), .op(n27591) );
  nand2_1 U31466 ( .ip1(n27592), .ip2(n27591), .op(n13450) );
endmodule

