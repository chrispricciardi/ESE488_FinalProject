
module mult ( clk, reset, in, w, out );
  input [15:0] in;
  input [15:0] w;
  output [15:0] out;
  input clk, reset;
  wire   \layer1[15][23] , \layer1[15][22] , \layer1[15][21] ,
         \layer1[15][20] , \layer1[15][19] , \layer1[15][18] ,
         \layer1[15][17] , \layer1[15][16] , \layer1[15][15] ,
         \layer1[14][23] , \layer1[14][22] , \layer1[14][21] ,
         \layer1[14][20] , \layer1[14][19] , \layer1[14][18] ,
         \layer1[14][17] , \layer1[14][16] , \layer1[14][15] ,
         \layer1[13][23] , \layer1[13][22] , \layer1[13][21] ,
         \layer1[13][20] , \layer1[13][19] , \layer1[13][18] ,
         \layer1[13][17] , \layer1[13][16] , \layer1[13][15] ,
         \layer1[13][14] , \layer1[13][13] , \layer1[12][23] ,
         \layer1[12][22] , \layer1[12][21] , \layer1[12][20] ,
         \layer1[12][19] , \layer1[12][18] , \layer1[12][17] ,
         \layer1[12][16] , \layer1[12][15] , \layer1[12][14] ,
         \layer1[12][13] , \layer1[11][23] , \layer1[11][22] ,
         \layer1[11][21] , \layer1[11][20] , \layer1[11][19] ,
         \layer1[11][18] , \layer1[11][17] , \layer1[11][16] ,
         \layer1[11][15] , \layer1[11][14] , \layer1[11][13] ,
         \layer1[11][12] , \layer1[11][11] , \layer1[10][23] ,
         \layer1[10][22] , \layer1[10][21] , \layer1[10][20] ,
         \layer1[10][19] , \layer1[10][18] , \layer1[10][17] ,
         \layer1[10][16] , \layer1[10][15] , \layer1[10][14] ,
         \layer1[10][13] , \layer1[10][12] , \layer1[10][11] , \layer1[9][23] ,
         \layer1[9][22] , \layer1[9][21] , \layer1[9][20] , \layer1[9][19] ,
         \layer1[9][18] , \layer1[9][17] , \layer1[9][16] , \layer1[9][15] ,
         \layer1[9][14] , \layer1[9][13] , \layer1[9][12] , \layer1[9][11] ,
         \layer1[9][10] , \layer1[9][9] , \layer1[8][23] , \layer1[8][22] ,
         \layer1[8][21] , \layer1[8][20] , \layer1[8][19] , \layer1[8][18] ,
         \layer1[8][17] , \layer1[8][16] , \layer1[8][15] , \layer1[8][14] ,
         \layer1[8][13] , \layer1[8][12] , \layer1[8][11] , \layer1[8][10] ,
         \layer1[8][9] , \layer1[7][22] , \layer1[7][21] , \layer1[7][20] ,
         \layer1[7][19] , \layer1[7][18] , \layer1[7][17] , \layer1[7][16] ,
         \layer1[7][15] , \layer1[7][14] , \layer1[7][13] , \layer1[7][12] ,
         \layer1[7][11] , \layer1[7][10] , \layer1[7][9] , \layer1[7][8] ,
         \layer1[7][7] , \layer1[6][21] , \layer1[6][20] , \layer1[6][19] ,
         \layer1[6][18] , \layer1[6][17] , \layer1[6][16] , \layer1[6][15] ,
         \layer1[6][14] , \layer1[6][13] , \layer1[6][12] , \layer1[6][11] ,
         \layer1[6][10] , \layer1[6][9] , \layer1[6][8] , \layer1[6][7] ,
         \layer1[5][20] , \layer1[5][19] , \layer1[5][18] , \layer1[5][17] ,
         \layer1[5][16] , \layer1[5][15] , \layer1[5][14] , \layer1[5][13] ,
         \layer1[5][12] , \layer1[5][11] , \layer1[5][10] , \layer1[5][9] ,
         \layer1[5][8] , \layer1[5][7] , \layer1[5][6] , \layer1[5][5] ,
         \layer1[4][19] , \layer1[4][18] , \layer1[4][17] , \layer1[4][16] ,
         \layer1[4][15] , \layer1[4][14] , \layer1[4][13] , \layer1[4][12] ,
         \layer1[4][11] , \layer1[4][10] , \layer1[4][9] , \layer1[4][8] ,
         \layer1[4][7] , \layer1[4][6] , \layer1[4][5] , \layer1[3][18] ,
         \layer1[3][17] , \layer1[3][16] , \layer1[3][15] , \layer1[3][14] ,
         \layer1[3][13] , \layer1[3][12] , \layer1[3][11] , \layer1[3][10] ,
         \layer1[3][9] , \layer1[3][8] , \layer1[3][7] , \layer1[3][6] ,
         \layer1[3][5] , \layer1[3][4] , \layer1[3][3] , \layer1[2][17] ,
         \layer1[2][16] , \layer1[2][15] , \layer1[2][14] , \layer1[2][13] ,
         \layer1[2][12] , \layer1[2][11] , \layer1[2][10] , \layer1[2][9] ,
         \layer1[2][8] , \layer1[2][7] , \layer1[2][6] , \layer1[2][5] ,
         \layer1[2][4] , \layer1[2][3] , \layer1[1][16] , \layer1[1][15] ,
         \layer1[1][14] , \layer1[1][13] , \layer1[1][12] , \layer1[1][11] ,
         \layer1[1][10] , \layer1[1][9] , \layer1[1][8] , \layer1[1][7] ,
         \layer1[1][6] , \layer1[1][5] , \layer1[1][4] , \layer1[1][3] ,
         \layer1[1][2] , \layer1[1][1] , \layer1[0][16] , \layer1[0][15] ,
         \layer1[0][14] , \layer1[0][13] , \layer1[0][12] , \layer1[0][11] ,
         \layer1[0][10] , \layer1[0][9] , \layer1[0][8] , \layer1[0][7] ,
         \layer1[0][6] , \layer1[0][5] , \layer1[0][4] , \layer1[0][3] ,
         \layer1[0][2] , \layer1[0][1] , N293, N327, N361, N395, N429, N463,
         N497, \layer2[7][23] , \layer2[7][22] , \layer2[7][21] ,
         \layer2[7][20] , \layer2[7][19] , \layer2[7][18] , \layer2[7][17] ,
         \layer2[7][16] , \layer2[7][15] , \layer2[7][14] , \layer2[6][23] ,
         \layer2[6][22] , \layer2[6][21] , \layer2[6][20] , \layer2[6][19] ,
         \layer2[6][18] , \layer2[6][17] , \layer2[6][16] , \layer2[6][15] ,
         \layer2[6][14] , \layer2[5][23] , \layer2[5][22] , \layer2[5][21] ,
         \layer2[5][20] , \layer2[5][19] , \layer2[5][18] , \layer2[5][17] ,
         \layer2[5][16] , \layer2[5][15] , \layer2[5][14] , \layer2[5][13] ,
         \layer2[5][12] , \layer2[5][11] , \layer2[5][10] , \layer2[4][23] ,
         \layer2[4][22] , \layer2[4][21] , \layer2[4][20] , \layer2[4][19] ,
         \layer2[4][18] , \layer2[4][17] , \layer2[4][16] , \layer2[4][15] ,
         \layer2[4][14] , \layer2[4][13] , \layer2[4][12] , \layer2[4][11] ,
         \layer2[4][10] , \layer2[3][23] , \layer2[3][22] , \layer2[3][21] ,
         \layer2[3][20] , \layer2[3][19] , \layer2[3][18] , \layer2[3][17] ,
         \layer2[3][16] , \layer2[3][15] , \layer2[3][14] , \layer2[3][13] ,
         \layer2[3][12] , \layer2[3][11] , \layer2[3][10] , \layer2[3][9] ,
         \layer2[3][8] , \layer2[3][7] , \layer2[3][6] , \layer2[2][21] ,
         \layer2[2][20] , \layer2[2][19] , \layer2[2][18] , \layer2[2][17] ,
         \layer2[2][16] , \layer2[2][15] , \layer2[2][14] , \layer2[2][13] ,
         \layer2[2][12] , \layer2[2][11] , \layer2[2][10] , \layer2[2][9] ,
         \layer2[2][8] , \layer2[2][7] , \layer2[2][6] , \layer2[1][19] ,
         \layer2[1][18] , \layer2[1][17] , \layer2[1][16] , \layer2[1][15] ,
         \layer2[1][14] , \layer2[1][13] , \layer2[1][12] , \layer2[1][11] ,
         \layer2[1][10] , \layer2[1][9] , \layer2[1][8] , \layer2[1][7] ,
         \layer2[1][6] , \layer2[1][5] , \layer2[1][4] , \layer2[1][3] ,
         \layer2[1][2] , \layer2[0][17] , \layer2[0][16] , \layer2[0][15] ,
         \layer2[0][14] , \layer2[0][13] , \layer2[0][12] , \layer2[0][11] ,
         \layer2[0][10] , \layer2[0][9] , \layer2[0][8] , \layer2[0][7] ,
         \layer2[0][6] , \layer2[0][5] , \layer2[0][4] , \layer2[0][3] ,
         \layer2[0][2] , N551, N552, N587, N588, N623, N624, \layer3[3][23] ,
         \layer3[3][22] , \layer3[3][21] , \layer3[3][20] , \layer3[3][19] ,
         \layer3[3][18] , \layer3[3][17] , \layer3[3][16] , \layer3[3][15] ,
         \layer3[3][14] , \layer3[3][13] , \layer3[3][12] , \layer3[2][23] ,
         \layer3[2][22] , \layer3[2][21] , \layer3[2][20] , \layer3[2][19] ,
         \layer3[2][18] , \layer3[2][17] , \layer3[2][16] , \layer3[2][15] ,
         \layer3[2][14] , \layer3[2][13] , \layer3[2][12] , \layer3[1][23] ,
         \layer3[1][22] , \layer3[1][21] , \layer3[1][20] , \layer3[1][19] ,
         \layer3[1][18] , \layer3[1][17] , \layer3[1][16] , \layer3[1][15] ,
         \layer3[1][14] , \layer3[1][13] , \layer3[1][12] , \layer3[1][11] ,
         \layer3[1][10] , \layer3[1][9] , \layer3[1][8] , \layer3[1][7] ,
         \layer3[1][6] , \layer3[1][5] , \layer3[1][4] , \layer3[0][20] ,
         \layer3[0][19] , \layer3[0][18] , \layer3[0][17] , \layer3[0][16] ,
         \layer3[0][15] , \layer3[0][14] , \layer3[0][13] , \layer3[0][12] ,
         \layer3[0][11] , \layer3[0][10] , \layer3[0][9] , \layer3[0][8] ,
         \layer3[0][7] , \layer3[0][6] , \layer3[0][5] , \layer3[0][4] , N675,
         N676, N677, N678, \layer4[1][23] , \layer4[1][22] , \layer4[1][21] ,
         \layer4[1][20] , \layer4[1][19] , \layer4[1][18] , \layer4[1][17] ,
         \layer4[1][16] , \layer4[1][15] , \layer4[1][14] , \layer4[1][13] ,
         \layer4[1][12] , \layer4[1][11] , \layer4[1][10] , \layer4[1][9] ,
         \layer4[1][8] , \layer4[0][23] , \layer4[0][22] , \layer4[0][21] ,
         \layer4[0][20] , \layer4[0][19] , \layer4[0][18] , \layer4[0][17] ,
         \layer4[0][16] , \layer4[0][15] , \layer4[0][14] , \layer4[0][13] ,
         \layer4[0][12] , \layer4[0][11] , \layer4[0][10] , \layer4[0][9] ,
         \layer4[0][8] , N707, N708, N709, N710, N711, N712, N713, N714, N715,
         N716, N717, N718, N719, N720, N721, N722, N724, N725, N726, N727,
         N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738,
         N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749,
         N750, N751, N752, N753, N754, N755, N756, N757, N758, N759, N760,
         N761, N762, N763, N764, N765, N766, N767, N768, N769, N770, N771,
         N772, N773, N774, N775, N776, N777, N778, N779, N780, N781, N782,
         N783, N784, N785, N786, N787, N788, N789, N790, N791, N792, N793,
         N794, N795, N796, N797, N798, N799, N800, N801, N802, N803, N804,
         N805, N806, N807, N808, N809, N810, N811, N812, N813, N814, N815,
         N816, N817, N818, N819, N820, N821, N822, N823, N824, N825, N826,
         N827, N828, N829, N830, N831, N832, N833, N834, N835, N836, N837,
         N838, N839, N840, N841, N842, N843, N844, N845, N846, N847, N848,
         N849, N850, N851, N852, N853, N854, N855, N856, N857, N858, N859,
         N860, N861, N862, N863, N864, N865, N866, N867, N868, N869, N870,
         N871, N872, N873, N874, N875, N876, N877, N878, N879, N880, N881,
         N883, N884, N885, N886, N887, N888, N889, N890, N891, N892, N893,
         N894, N895, N896, N899, N900, N901, N902, N903, N904, N905, N906,
         N907, N908, N909, N910, N911, N915, N916, N917, N918, N919, N920,
         N921, N922, N923, N924, N925, N926, N931, N932, N933, N934, N935,
         N936, N937, N938, N939, N940, N941, N947, N948, N949, N950, N951,
         N952, N953, N954, N955, N956, N963, N964, N965, N966, N967, N968,
         N969, N970, N971, N981, N982, N983, N984, N985, N986, N987, N988,
         N989, N990, N991, N992, N993, N994, N995, N996, N1013, N1014, N1015,
         N1016, N1017, N1018, N1019, N1020, N1021, N1022, N1023, N1024, N1025,
         N1026, N1027, N1028, N1029, N1030, N1047, N1048, N1049, N1050, N1051,
         N1052, N1053, N1054, N1055, N1056, N1057, N1058, N1059, N1060, N1061,
         N1062, N1063, N1064, N1081, N1082, N1083, N1084, N1085, N1086, N1087,
         N1088, N1089, N1090, N1091, N1092, N1093, N1094, N1095, N1096, N1097,
         N1098, N1115, N1116, N1117, N1118, N1119, N1120, N1121, N1122, N1123,
         N1124, N1125, N1126, N1127, N1128, N1129, N1130, N1149, N1150, N1151,
         N1152, N1153, N1154, N1155, N1156, N1157, N1158, N1159, N1160, N1161,
         N1162, N1183, N1184, N1185, N1186, N1187, N1188, N1189, N1190, N1191,
         N1192, N1193, N1194, N1217, N1218, N1219, N1220, N1221, N1222, N1223,
         N1224, N1225, N1226, N1239, N1240, N1241, N1242, N1243, N1244, N1245,
         N1246, N1247, N1248, N1249, N1250, N1251, N1252, N1253, N1254, N1255,
         N1271, N1272, N1273, N1274, N1275, N1276, N1277, N1278, N1279, N1280,
         N1281, N1282, N1283, N1284, N1285, N1286, N1287, N1288, N1289, N1290,
         N1307, N1308, N1309, N1310, N1311, N1312, N1313, N1314, N1315, N1316,
         N1317, N1318, N1319, N1320, N1321, N1322, N1343, N1344, N1345, N1346,
         N1347, N1348, N1349, N1350, N1351, N1352, N1353, N1354, N1371, N1372,
         N1373, N1374, N1375, N1376, N1377, N1378, N1379, N1380, N1381, N1382,
         N1383, N1384, N1385, N1386, N1395, N1396, N1397, N1398, N1399, N1400,
         N1401, N1402, N1403, N1404, N1405, N1406, N1407, N1408, N1409, N1410,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840;

  dp_1 \layer5_reg[23]  ( .ip(N722), .ck(clk), .q(out[15]) );
  dp_1 \layer5_reg[22]  ( .ip(N721), .ck(clk), .q(out[14]) );
  dp_1 \layer5_reg[21]  ( .ip(N720), .ck(clk), .q(out[13]) );
  dp_1 \layer5_reg[20]  ( .ip(N719), .ck(clk), .q(out[12]) );
  dp_1 \layer5_reg[19]  ( .ip(N718), .ck(clk), .q(out[11]) );
  dp_1 \layer5_reg[18]  ( .ip(N717), .ck(clk), .q(out[10]) );
  dp_1 \layer5_reg[17]  ( .ip(N716), .ck(clk), .q(out[9]) );
  dp_1 \layer5_reg[16]  ( .ip(N715), .ck(clk), .q(out[8]) );
  dp_1 \layer5_reg[15]  ( .ip(N714), .ck(clk), .q(out[7]) );
  dp_1 \layer5_reg[14]  ( .ip(N713), .ck(clk), .q(out[6]) );
  dp_1 \layer5_reg[13]  ( .ip(N712), .ck(clk), .q(out[5]) );
  dp_1 \layer5_reg[12]  ( .ip(N711), .ck(clk), .q(out[4]) );
  dp_1 \layer5_reg[11]  ( .ip(N710), .ck(clk), .q(out[3]) );
  dp_1 \layer5_reg[10]  ( .ip(N709), .ck(clk), .q(out[2]) );
  dp_1 \layer5_reg[9]  ( .ip(N708), .ck(clk), .q(out[1]) );
  dp_1 \layer5_reg[8]  ( .ip(N707), .ck(clk), .q(out[0]) );
  dp_1 \layer4_reg[1][23]  ( .ip(N1410), .ck(clk), .q(\layer4[1][23] ) );
  dp_1 \layer4_reg[1][22]  ( .ip(N1409), .ck(clk), .q(\layer4[1][22] ) );
  dp_1 \layer4_reg[1][21]  ( .ip(N1408), .ck(clk), .q(\layer4[1][21] ) );
  dp_1 \layer4_reg[1][20]  ( .ip(N1407), .ck(clk), .q(\layer4[1][20] ) );
  dp_1 \layer4_reg[1][19]  ( .ip(N1406), .ck(clk), .q(\layer4[1][19] ) );
  dp_1 \layer4_reg[1][18]  ( .ip(N1405), .ck(clk), .q(\layer4[1][18] ) );
  dp_1 \layer4_reg[1][17]  ( .ip(N1404), .ck(clk), .q(\layer4[1][17] ) );
  dp_1 \layer4_reg[1][16]  ( .ip(N1403), .ck(clk), .q(\layer4[1][16] ) );
  dp_1 \layer4_reg[1][15]  ( .ip(N1402), .ck(clk), .q(\layer4[1][15] ) );
  dp_1 \layer4_reg[1][14]  ( .ip(N1401), .ck(clk), .q(\layer4[1][14] ) );
  dp_1 \layer4_reg[1][13]  ( .ip(N1400), .ck(clk), .q(\layer4[1][13] ) );
  dp_1 \layer4_reg[1][12]  ( .ip(N1399), .ck(clk), .q(\layer4[1][12] ) );
  dp_1 \layer4_reg[1][11]  ( .ip(N1398), .ck(clk), .q(\layer4[1][11] ) );
  dp_1 \layer4_reg[1][10]  ( .ip(N1397), .ck(clk), .q(\layer4[1][10] ) );
  dp_1 \layer4_reg[1][9]  ( .ip(N1396), .ck(clk), .q(\layer4[1][9] ) );
  dp_1 \layer4_reg[1][8]  ( .ip(N1395), .ck(clk), .q(\layer4[1][8] ) );
  dp_1 \layer4_reg[0][23]  ( .ip(N1386), .ck(clk), .q(\layer4[0][23] ) );
  dp_1 \layer4_reg[0][22]  ( .ip(N1385), .ck(clk), .q(\layer4[0][22] ) );
  dp_1 \layer4_reg[0][21]  ( .ip(N1384), .ck(clk), .q(\layer4[0][21] ) );
  dp_1 \layer4_reg[0][20]  ( .ip(N1383), .ck(clk), .q(\layer4[0][20] ) );
  dp_1 \layer4_reg[0][19]  ( .ip(N1382), .ck(clk), .q(\layer4[0][19] ) );
  dp_1 \layer4_reg[0][18]  ( .ip(N1381), .ck(clk), .q(\layer4[0][18] ) );
  dp_1 \layer4_reg[0][17]  ( .ip(N1380), .ck(clk), .q(\layer4[0][17] ) );
  dp_1 \layer4_reg[0][16]  ( .ip(N1379), .ck(clk), .q(\layer4[0][16] ) );
  dp_1 \layer4_reg[0][15]  ( .ip(N1378), .ck(clk), .q(\layer4[0][15] ) );
  dp_1 \layer4_reg[0][14]  ( .ip(N1377), .ck(clk), .q(\layer4[0][14] ) );
  dp_1 \layer4_reg[0][13]  ( .ip(N1376), .ck(clk), .q(\layer4[0][13] ) );
  dp_1 \layer4_reg[0][12]  ( .ip(N1375), .ck(clk), .q(\layer4[0][12] ) );
  dp_1 \layer4_reg[0][11]  ( .ip(N1374), .ck(clk), .q(\layer4[0][11] ) );
  dp_1 \layer4_reg[0][10]  ( .ip(N1373), .ck(clk), .q(\layer4[0][10] ) );
  dp_1 \layer4_reg[0][9]  ( .ip(N1372), .ck(clk), .q(\layer4[0][9] ) );
  dp_1 \layer4_reg[0][8]  ( .ip(N1371), .ck(clk), .q(\layer4[0][8] ) );
  dp_1 \layer2_reg[7][23]  ( .ip(N1226), .ck(clk), .q(\layer2[7][23] ) );
  dp_1 \layer2_reg[7][22]  ( .ip(N1225), .ck(clk), .q(\layer2[7][22] ) );
  dp_1 \layer2_reg[7][21]  ( .ip(N1224), .ck(clk), .q(\layer2[7][21] ) );
  dp_1 \layer2_reg[7][20]  ( .ip(N1223), .ck(clk), .q(\layer2[7][20] ) );
  dp_1 \layer2_reg[7][19]  ( .ip(N1222), .ck(clk), .q(\layer2[7][19] ) );
  dp_1 \layer2_reg[7][18]  ( .ip(N1221), .ck(clk), .q(\layer2[7][18] ) );
  dp_1 \layer2_reg[7][17]  ( .ip(N1220), .ck(clk), .q(\layer2[7][17] ) );
  dp_1 \layer2_reg[7][16]  ( .ip(N1219), .ck(clk), .q(\layer2[7][16] ) );
  dp_1 \layer2_reg[7][15]  ( .ip(N1218), .ck(clk), .q(\layer2[7][15] ) );
  dp_1 \layer2_reg[7][14]  ( .ip(N1217), .ck(clk), .q(\layer2[7][14] ) );
  dp_1 \layer2_reg[6][23]  ( .ip(N1194), .ck(clk), .q(\layer2[6][23] ) );
  dp_1 \layer2_reg[6][22]  ( .ip(N1193), .ck(clk), .q(\layer2[6][22] ) );
  dp_1 \layer2_reg[6][21]  ( .ip(N1192), .ck(clk), .q(\layer2[6][21] ) );
  dp_1 \layer2_reg[6][20]  ( .ip(N1191), .ck(clk), .q(\layer2[6][20] ) );
  dp_1 \layer2_reg[6][19]  ( .ip(N1190), .ck(clk), .q(\layer2[6][19] ) );
  dp_1 \layer2_reg[6][18]  ( .ip(N1189), .ck(clk), .q(\layer2[6][18] ) );
  dp_1 \layer2_reg[6][17]  ( .ip(N1188), .ck(clk), .q(\layer2[6][17] ) );
  dp_1 \layer2_reg[6][16]  ( .ip(N1187), .ck(clk), .q(\layer2[6][16] ) );
  dp_1 \layer2_reg[6][15]  ( .ip(N1186), .ck(clk), .q(\layer2[6][15] ) );
  dp_1 \layer2_reg[6][14]  ( .ip(N1185), .ck(clk), .q(\layer2[6][14] ) );
  dp_1 \layer2_reg[6][13]  ( .ip(N1184), .ck(clk), .q(N624) );
  dp_1 \layer2_reg[6][12]  ( .ip(N1183), .ck(clk), .q(N623) );
  dp_1 \layer2_reg[5][23]  ( .ip(N1162), .ck(clk), .q(\layer2[5][23] ) );
  dp_1 \layer2_reg[5][22]  ( .ip(N1161), .ck(clk), .q(\layer2[5][22] ) );
  dp_1 \layer2_reg[5][21]  ( .ip(N1160), .ck(clk), .q(\layer2[5][21] ) );
  dp_1 \layer2_reg[5][20]  ( .ip(N1159), .ck(clk), .q(\layer2[5][20] ) );
  dp_1 \layer2_reg[5][19]  ( .ip(N1158), .ck(clk), .q(\layer2[5][19] ) );
  dp_1 \layer2_reg[5][18]  ( .ip(N1157), .ck(clk), .q(\layer2[5][18] ) );
  dp_1 \layer2_reg[5][17]  ( .ip(N1156), .ck(clk), .q(\layer2[5][17] ) );
  dp_1 \layer2_reg[5][16]  ( .ip(N1155), .ck(clk), .q(\layer2[5][16] ) );
  dp_1 \layer2_reg[5][15]  ( .ip(N1154), .ck(clk), .q(\layer2[5][15] ) );
  dp_1 \layer2_reg[5][14]  ( .ip(N1153), .ck(clk), .q(\layer2[5][14] ) );
  dp_1 \layer2_reg[5][13]  ( .ip(N1152), .ck(clk), .q(\layer2[5][13] ) );
  dp_1 \layer2_reg[5][12]  ( .ip(N1151), .ck(clk), .q(\layer2[5][12] ) );
  dp_1 \layer2_reg[5][11]  ( .ip(N1150), .ck(clk), .q(\layer2[5][11] ) );
  dp_1 \layer2_reg[5][10]  ( .ip(N1149), .ck(clk), .q(\layer2[5][10] ) );
  dp_1 \layer2_reg[4][23]  ( .ip(N1130), .ck(clk), .q(\layer2[4][23] ) );
  dp_1 \layer2_reg[4][22]  ( .ip(N1129), .ck(clk), .q(\layer2[4][22] ) );
  dp_1 \layer2_reg[4][21]  ( .ip(N1128), .ck(clk), .q(\layer2[4][21] ) );
  dp_1 \layer2_reg[4][20]  ( .ip(N1127), .ck(clk), .q(\layer2[4][20] ) );
  dp_1 \layer2_reg[4][19]  ( .ip(N1126), .ck(clk), .q(\layer2[4][19] ) );
  dp_1 \layer2_reg[4][18]  ( .ip(N1125), .ck(clk), .q(\layer2[4][18] ) );
  dp_1 \layer2_reg[4][17]  ( .ip(N1124), .ck(clk), .q(\layer2[4][17] ) );
  dp_1 \layer2_reg[4][16]  ( .ip(N1123), .ck(clk), .q(\layer2[4][16] ) );
  dp_1 \layer2_reg[4][15]  ( .ip(N1122), .ck(clk), .q(\layer2[4][15] ) );
  dp_1 \layer2_reg[4][14]  ( .ip(N1121), .ck(clk), .q(\layer2[4][14] ) );
  dp_1 \layer2_reg[4][13]  ( .ip(N1120), .ck(clk), .q(\layer2[4][13] ) );
  dp_1 \layer2_reg[4][12]  ( .ip(N1119), .ck(clk), .q(\layer2[4][12] ) );
  dp_1 \layer2_reg[4][11]  ( .ip(N1118), .ck(clk), .q(\layer2[4][11] ) );
  dp_1 \layer2_reg[4][10]  ( .ip(N1117), .ck(clk), .q(\layer2[4][10] ) );
  dp_1 \layer2_reg[4][9]  ( .ip(N1116), .ck(clk), .q(N588) );
  dp_1 \layer2_reg[4][8]  ( .ip(N1115), .ck(clk), .q(N587) );
  dp_1 \layer2_reg[3][23]  ( .ip(N1098), .ck(clk), .q(\layer2[3][23] ) );
  dp_1 \layer2_reg[3][22]  ( .ip(N1097), .ck(clk), .q(\layer2[3][22] ) );
  dp_1 \layer2_reg[3][21]  ( .ip(N1096), .ck(clk), .q(\layer2[3][21] ) );
  dp_1 \layer2_reg[3][20]  ( .ip(N1095), .ck(clk), .q(\layer2[3][20] ) );
  dp_1 \layer2_reg[3][19]  ( .ip(N1094), .ck(clk), .q(\layer2[3][19] ) );
  dp_1 \layer2_reg[3][18]  ( .ip(N1093), .ck(clk), .q(\layer2[3][18] ) );
  dp_1 \layer2_reg[3][17]  ( .ip(N1092), .ck(clk), .q(\layer2[3][17] ) );
  dp_1 \layer2_reg[3][16]  ( .ip(N1091), .ck(clk), .q(\layer2[3][16] ) );
  dp_1 \layer2_reg[3][15]  ( .ip(N1090), .ck(clk), .q(\layer2[3][15] ) );
  dp_1 \layer2_reg[3][14]  ( .ip(N1089), .ck(clk), .q(\layer2[3][14] ) );
  dp_1 \layer2_reg[3][13]  ( .ip(N1088), .ck(clk), .q(\layer2[3][13] ) );
  dp_1 \layer2_reg[3][12]  ( .ip(N1087), .ck(clk), .q(\layer2[3][12] ) );
  dp_1 \layer2_reg[3][11]  ( .ip(N1086), .ck(clk), .q(\layer2[3][11] ) );
  dp_1 \layer2_reg[3][10]  ( .ip(N1085), .ck(clk), .q(\layer2[3][10] ) );
  dp_1 \layer2_reg[3][9]  ( .ip(N1084), .ck(clk), .q(\layer2[3][9] ) );
  dp_1 \layer2_reg[3][8]  ( .ip(N1083), .ck(clk), .q(\layer2[3][8] ) );
  dp_1 \layer2_reg[3][7]  ( .ip(N1082), .ck(clk), .q(\layer2[3][7] ) );
  dp_1 \layer2_reg[3][6]  ( .ip(N1081), .ck(clk), .q(\layer2[3][6] ) );
  dp_1 \layer2_reg[2][21]  ( .ip(N1064), .ck(clk), .q(\layer2[2][21] ) );
  dp_1 \layer2_reg[2][20]  ( .ip(N1063), .ck(clk), .q(\layer2[2][20] ) );
  dp_1 \layer2_reg[2][19]  ( .ip(N1062), .ck(clk), .q(\layer2[2][19] ) );
  dp_1 \layer2_reg[2][18]  ( .ip(N1061), .ck(clk), .q(\layer2[2][18] ) );
  dp_1 \layer2_reg[2][17]  ( .ip(N1060), .ck(clk), .q(\layer2[2][17] ) );
  dp_1 \layer2_reg[2][16]  ( .ip(N1059), .ck(clk), .q(\layer2[2][16] ) );
  dp_1 \layer2_reg[2][15]  ( .ip(N1058), .ck(clk), .q(\layer2[2][15] ) );
  dp_1 \layer2_reg[2][14]  ( .ip(N1057), .ck(clk), .q(\layer2[2][14] ) );
  dp_1 \layer2_reg[2][13]  ( .ip(N1056), .ck(clk), .q(\layer2[2][13] ) );
  dp_1 \layer2_reg[2][12]  ( .ip(N1055), .ck(clk), .q(\layer2[2][12] ) );
  dp_1 \layer2_reg[2][11]  ( .ip(N1054), .ck(clk), .q(\layer2[2][11] ) );
  dp_1 \layer2_reg[2][10]  ( .ip(N1053), .ck(clk), .q(\layer2[2][10] ) );
  dp_1 \layer2_reg[2][9]  ( .ip(N1052), .ck(clk), .q(\layer2[2][9] ) );
  dp_1 \layer2_reg[2][8]  ( .ip(N1051), .ck(clk), .q(\layer2[2][8] ) );
  dp_1 \layer2_reg[2][7]  ( .ip(N1050), .ck(clk), .q(\layer2[2][7] ) );
  dp_1 \layer2_reg[2][6]  ( .ip(N1049), .ck(clk), .q(\layer2[2][6] ) );
  dp_1 \layer2_reg[2][5]  ( .ip(N1048), .ck(clk), .q(N552) );
  dp_1 \layer2_reg[2][4]  ( .ip(N1047), .ck(clk), .q(N551) );
  dp_1 \layer2_reg[1][19]  ( .ip(N1030), .ck(clk), .q(\layer2[1][19] ) );
  dp_1 \layer2_reg[1][18]  ( .ip(N1029), .ck(clk), .q(\layer2[1][18] ) );
  dp_1 \layer2_reg[1][17]  ( .ip(N1028), .ck(clk), .q(\layer2[1][17] ) );
  dp_1 \layer2_reg[1][16]  ( .ip(N1027), .ck(clk), .q(\layer2[1][16] ) );
  dp_1 \layer2_reg[1][15]  ( .ip(N1026), .ck(clk), .q(\layer2[1][15] ) );
  dp_1 \layer2_reg[1][14]  ( .ip(N1025), .ck(clk), .q(\layer2[1][14] ) );
  dp_1 \layer2_reg[1][13]  ( .ip(N1024), .ck(clk), .q(\layer2[1][13] ) );
  dp_1 \layer2_reg[1][12]  ( .ip(N1023), .ck(clk), .q(\layer2[1][12] ) );
  dp_1 \layer2_reg[1][11]  ( .ip(N1022), .ck(clk), .q(\layer2[1][11] ) );
  dp_1 \layer2_reg[1][10]  ( .ip(N1021), .ck(clk), .q(\layer2[1][10] ) );
  dp_1 \layer2_reg[1][9]  ( .ip(N1020), .ck(clk), .q(\layer2[1][9] ) );
  dp_1 \layer2_reg[1][8]  ( .ip(N1019), .ck(clk), .q(\layer2[1][8] ) );
  dp_1 \layer2_reg[1][7]  ( .ip(N1018), .ck(clk), .q(\layer2[1][7] ) );
  dp_1 \layer2_reg[1][6]  ( .ip(N1017), .ck(clk), .q(\layer2[1][6] ) );
  dp_1 \layer2_reg[1][5]  ( .ip(N1016), .ck(clk), .q(\layer2[1][5] ) );
  dp_1 \layer2_reg[1][4]  ( .ip(N1015), .ck(clk), .q(\layer2[1][4] ) );
  dp_1 \layer2_reg[1][3]  ( .ip(N1014), .ck(clk), .q(\layer2[1][3] ) );
  dp_1 \layer2_reg[1][2]  ( .ip(N1013), .ck(clk), .q(\layer2[1][2] ) );
  dp_1 \layer2_reg[0][17]  ( .ip(N996), .ck(clk), .q(\layer2[0][17] ) );
  dp_1 \layer2_reg[0][16]  ( .ip(N995), .ck(clk), .q(\layer2[0][16] ) );
  dp_1 \layer2_reg[0][15]  ( .ip(N994), .ck(clk), .q(\layer2[0][15] ) );
  dp_1 \layer2_reg[0][14]  ( .ip(N993), .ck(clk), .q(\layer2[0][14] ) );
  dp_1 \layer2_reg[0][13]  ( .ip(N992), .ck(clk), .q(\layer2[0][13] ) );
  dp_1 \layer2_reg[0][12]  ( .ip(N991), .ck(clk), .q(\layer2[0][12] ) );
  dp_1 \layer2_reg[0][11]  ( .ip(N990), .ck(clk), .q(\layer2[0][11] ) );
  dp_1 \layer2_reg[0][10]  ( .ip(N989), .ck(clk), .q(\layer2[0][10] ) );
  dp_1 \layer2_reg[0][9]  ( .ip(N988), .ck(clk), .q(\layer2[0][9] ) );
  dp_1 \layer2_reg[0][8]  ( .ip(N987), .ck(clk), .q(\layer2[0][8] ) );
  dp_1 \layer2_reg[0][7]  ( .ip(N986), .ck(clk), .q(\layer2[0][7] ) );
  dp_1 \layer2_reg[0][6]  ( .ip(N985), .ck(clk), .q(\layer2[0][6] ) );
  dp_1 \layer2_reg[0][5]  ( .ip(N984), .ck(clk), .q(\layer2[0][5] ) );
  dp_1 \layer2_reg[0][4]  ( .ip(N983), .ck(clk), .q(\layer2[0][4] ) );
  dp_1 \layer2_reg[0][3]  ( .ip(N982), .ck(clk), .q(\layer2[0][3] ) );
  dp_1 \layer2_reg[0][2]  ( .ip(N981), .ck(clk), .q(\layer2[0][2] ) );
  dp_1 \layer3_reg[3][23]  ( .ip(N1354), .ck(clk), .q(\layer3[3][23] ) );
  dp_1 \layer3_reg[3][22]  ( .ip(N1353), .ck(clk), .q(\layer3[3][22] ) );
  dp_1 \layer3_reg[3][21]  ( .ip(N1352), .ck(clk), .q(\layer3[3][21] ) );
  dp_1 \layer3_reg[3][20]  ( .ip(N1351), .ck(clk), .q(\layer3[3][20] ) );
  dp_1 \layer3_reg[3][19]  ( .ip(N1350), .ck(clk), .q(\layer3[3][19] ) );
  dp_1 \layer3_reg[3][18]  ( .ip(N1349), .ck(clk), .q(\layer3[3][18] ) );
  dp_1 \layer3_reg[3][17]  ( .ip(N1348), .ck(clk), .q(\layer3[3][17] ) );
  dp_1 \layer3_reg[3][16]  ( .ip(N1347), .ck(clk), .q(\layer3[3][16] ) );
  dp_1 \layer3_reg[3][15]  ( .ip(N1346), .ck(clk), .q(\layer3[3][15] ) );
  dp_1 \layer3_reg[3][14]  ( .ip(N1345), .ck(clk), .q(\layer3[3][14] ) );
  dp_1 \layer3_reg[3][13]  ( .ip(N1344), .ck(clk), .q(\layer3[3][13] ) );
  dp_1 \layer3_reg[3][12]  ( .ip(N1343), .ck(clk), .q(\layer3[3][12] ) );
  dp_1 \layer3_reg[2][23]  ( .ip(N1322), .ck(clk), .q(\layer3[2][23] ) );
  dp_1 \layer3_reg[2][22]  ( .ip(N1321), .ck(clk), .q(\layer3[2][22] ) );
  dp_1 \layer3_reg[2][21]  ( .ip(N1320), .ck(clk), .q(\layer3[2][21] ) );
  dp_1 \layer3_reg[2][20]  ( .ip(N1319), .ck(clk), .q(\layer3[2][20] ) );
  dp_1 \layer3_reg[2][19]  ( .ip(N1318), .ck(clk), .q(\layer3[2][19] ) );
  dp_1 \layer3_reg[2][18]  ( .ip(N1317), .ck(clk), .q(\layer3[2][18] ) );
  dp_1 \layer3_reg[2][17]  ( .ip(N1316), .ck(clk), .q(\layer3[2][17] ) );
  dp_1 \layer3_reg[2][16]  ( .ip(N1315), .ck(clk), .q(\layer3[2][16] ) );
  dp_1 \layer3_reg[2][15]  ( .ip(N1314), .ck(clk), .q(\layer3[2][15] ) );
  dp_1 \layer3_reg[2][14]  ( .ip(N1313), .ck(clk), .q(\layer3[2][14] ) );
  dp_1 \layer3_reg[2][13]  ( .ip(N1312), .ck(clk), .q(\layer3[2][13] ) );
  dp_1 \layer3_reg[2][12]  ( .ip(N1311), .ck(clk), .q(\layer3[2][12] ) );
  dp_1 \layer3_reg[2][11]  ( .ip(N1310), .ck(clk), .q(N678) );
  dp_1 \layer3_reg[2][10]  ( .ip(N1309), .ck(clk), .q(N677) );
  dp_1 \layer3_reg[2][9]  ( .ip(N1308), .ck(clk), .q(N676) );
  dp_1 \layer3_reg[2][8]  ( .ip(N1307), .ck(clk), .q(N675) );
  dp_1 \layer3_reg[1][23]  ( .ip(N1290), .ck(clk), .q(\layer3[1][23] ) );
  dp_1 \layer3_reg[1][22]  ( .ip(N1289), .ck(clk), .q(\layer3[1][22] ) );
  dp_1 \layer3_reg[1][21]  ( .ip(N1288), .ck(clk), .q(\layer3[1][21] ) );
  dp_1 \layer3_reg[1][20]  ( .ip(N1287), .ck(clk), .q(\layer3[1][20] ) );
  dp_1 \layer3_reg[1][19]  ( .ip(N1286), .ck(clk), .q(\layer3[1][19] ) );
  dp_1 \layer3_reg[1][18]  ( .ip(N1285), .ck(clk), .q(\layer3[1][18] ) );
  dp_1 \layer3_reg[1][17]  ( .ip(N1284), .ck(clk), .q(\layer3[1][17] ) );
  dp_1 \layer3_reg[1][16]  ( .ip(N1283), .ck(clk), .q(\layer3[1][16] ) );
  dp_1 \layer3_reg[1][15]  ( .ip(N1282), .ck(clk), .q(\layer3[1][15] ) );
  dp_1 \layer3_reg[1][14]  ( .ip(N1281), .ck(clk), .q(\layer3[1][14] ) );
  dp_1 \layer3_reg[1][13]  ( .ip(N1280), .ck(clk), .q(\layer3[1][13] ) );
  dp_1 \layer3_reg[1][12]  ( .ip(N1279), .ck(clk), .q(\layer3[1][12] ) );
  dp_1 \layer3_reg[1][11]  ( .ip(N1278), .ck(clk), .q(\layer3[1][11] ) );
  dp_1 \layer3_reg[1][10]  ( .ip(N1277), .ck(clk), .q(\layer3[1][10] ) );
  dp_1 \layer3_reg[1][9]  ( .ip(N1276), .ck(clk), .q(\layer3[1][9] ) );
  dp_1 \layer3_reg[1][8]  ( .ip(N1275), .ck(clk), .q(\layer3[1][8] ) );
  dp_1 \layer3_reg[1][7]  ( .ip(N1274), .ck(clk), .q(\layer3[1][7] ) );
  dp_1 \layer3_reg[1][6]  ( .ip(N1273), .ck(clk), .q(\layer3[1][6] ) );
  dp_1 \layer3_reg[1][5]  ( .ip(N1272), .ck(clk), .q(\layer3[1][5] ) );
  dp_1 \layer3_reg[1][4]  ( .ip(N1271), .ck(clk), .q(\layer3[1][4] ) );
  dp_1 \layer3_reg[0][20]  ( .ip(N1255), .ck(clk), .q(\layer3[0][20] ) );
  dp_1 \layer3_reg[0][19]  ( .ip(N1254), .ck(clk), .q(\layer3[0][19] ) );
  dp_1 \layer3_reg[0][18]  ( .ip(N1253), .ck(clk), .q(\layer3[0][18] ) );
  dp_1 \layer3_reg[0][17]  ( .ip(N1252), .ck(clk), .q(\layer3[0][17] ) );
  dp_1 \layer3_reg[0][16]  ( .ip(N1251), .ck(clk), .q(\layer3[0][16] ) );
  dp_1 \layer3_reg[0][15]  ( .ip(N1250), .ck(clk), .q(\layer3[0][15] ) );
  dp_1 \layer3_reg[0][14]  ( .ip(N1249), .ck(clk), .q(\layer3[0][14] ) );
  dp_1 \layer3_reg[0][13]  ( .ip(N1248), .ck(clk), .q(\layer3[0][13] ) );
  dp_1 \layer3_reg[0][12]  ( .ip(N1247), .ck(clk), .q(\layer3[0][12] ) );
  dp_1 \layer3_reg[0][11]  ( .ip(N1246), .ck(clk), .q(\layer3[0][11] ) );
  dp_1 \layer3_reg[0][10]  ( .ip(N1245), .ck(clk), .q(\layer3[0][10] ) );
  dp_1 \layer3_reg[0][9]  ( .ip(N1244), .ck(clk), .q(\layer3[0][9] ) );
  dp_1 \layer3_reg[0][8]  ( .ip(N1243), .ck(clk), .q(\layer3[0][8] ) );
  dp_1 \layer3_reg[0][7]  ( .ip(N1242), .ck(clk), .q(\layer3[0][7] ) );
  dp_1 \layer3_reg[0][6]  ( .ip(N1241), .ck(clk), .q(\layer3[0][6] ) );
  dp_1 \layer3_reg[0][5]  ( .ip(N1240), .ck(clk), .q(\layer3[0][5] ) );
  dp_1 \layer3_reg[0][4]  ( .ip(N1239), .ck(clk), .q(\layer3[0][4] ) );
  dp_1 \layer1_reg[15][23]  ( .ip(N971), .ck(clk), .q(\layer1[15][23] ) );
  dp_1 \layer1_reg[15][22]  ( .ip(N970), .ck(clk), .q(\layer1[15][22] ) );
  dp_1 \layer1_reg[15][21]  ( .ip(N969), .ck(clk), .q(\layer1[15][21] ) );
  dp_1 \layer1_reg[15][20]  ( .ip(N968), .ck(clk), .q(\layer1[15][20] ) );
  dp_1 \layer1_reg[15][19]  ( .ip(N967), .ck(clk), .q(\layer1[15][19] ) );
  dp_1 \layer1_reg[15][18]  ( .ip(N966), .ck(clk), .q(\layer1[15][18] ) );
  dp_1 \layer1_reg[15][17]  ( .ip(N965), .ck(clk), .q(\layer1[15][17] ) );
  dp_1 \layer1_reg[15][16]  ( .ip(N964), .ck(clk), .q(\layer1[15][16] ) );
  dp_1 \layer1_reg[15][15]  ( .ip(N963), .ck(clk), .q(\layer1[15][15] ) );
  dp_1 \layer1_reg[14][23]  ( .ip(N956), .ck(clk), .q(\layer1[14][23] ) );
  dp_1 \layer1_reg[14][22]  ( .ip(N955), .ck(clk), .q(\layer1[14][22] ) );
  dp_1 \layer1_reg[14][21]  ( .ip(N954), .ck(clk), .q(\layer1[14][21] ) );
  dp_1 \layer1_reg[14][20]  ( .ip(N953), .ck(clk), .q(\layer1[14][20] ) );
  dp_1 \layer1_reg[14][19]  ( .ip(N952), .ck(clk), .q(\layer1[14][19] ) );
  dp_1 \layer1_reg[14][18]  ( .ip(N951), .ck(clk), .q(\layer1[14][18] ) );
  dp_1 \layer1_reg[14][17]  ( .ip(N950), .ck(clk), .q(\layer1[14][17] ) );
  dp_1 \layer1_reg[14][16]  ( .ip(N949), .ck(clk), .q(\layer1[14][16] ) );
  dp_1 \layer1_reg[14][15]  ( .ip(N948), .ck(clk), .q(\layer1[14][15] ) );
  dp_1 \layer1_reg[14][14]  ( .ip(N947), .ck(clk), .q(N497) );
  dp_1 \layer1_reg[13][23]  ( .ip(N941), .ck(clk), .q(\layer1[13][23] ) );
  dp_1 \layer1_reg[13][22]  ( .ip(N940), .ck(clk), .q(\layer1[13][22] ) );
  dp_1 \layer1_reg[13][21]  ( .ip(N939), .ck(clk), .q(\layer1[13][21] ) );
  dp_1 \layer1_reg[13][20]  ( .ip(N938), .ck(clk), .q(\layer1[13][20] ) );
  dp_1 \layer1_reg[13][19]  ( .ip(N937), .ck(clk), .q(\layer1[13][19] ) );
  dp_1 \layer1_reg[13][18]  ( .ip(N936), .ck(clk), .q(\layer1[13][18] ) );
  dp_1 \layer1_reg[13][17]  ( .ip(N935), .ck(clk), .q(\layer1[13][17] ) );
  dp_1 \layer1_reg[13][16]  ( .ip(N934), .ck(clk), .q(\layer1[13][16] ) );
  dp_1 \layer1_reg[13][15]  ( .ip(N933), .ck(clk), .q(\layer1[13][15] ) );
  dp_1 \layer1_reg[13][14]  ( .ip(N932), .ck(clk), .q(\layer1[13][14] ) );
  dp_1 \layer1_reg[13][13]  ( .ip(N931), .ck(clk), .q(\layer1[13][13] ) );
  dp_1 \layer1_reg[12][23]  ( .ip(N926), .ck(clk), .q(\layer1[12][23] ) );
  dp_1 \layer1_reg[12][22]  ( .ip(N925), .ck(clk), .q(\layer1[12][22] ) );
  dp_1 \layer1_reg[12][21]  ( .ip(N924), .ck(clk), .q(\layer1[12][21] ) );
  dp_1 \layer1_reg[12][20]  ( .ip(N923), .ck(clk), .q(\layer1[12][20] ) );
  dp_1 \layer1_reg[12][19]  ( .ip(N922), .ck(clk), .q(\layer1[12][19] ) );
  dp_1 \layer1_reg[12][18]  ( .ip(N921), .ck(clk), .q(\layer1[12][18] ) );
  dp_1 \layer1_reg[12][17]  ( .ip(N920), .ck(clk), .q(\layer1[12][17] ) );
  dp_1 \layer1_reg[12][16]  ( .ip(N919), .ck(clk), .q(\layer1[12][16] ) );
  dp_1 \layer1_reg[12][15]  ( .ip(N918), .ck(clk), .q(\layer1[12][15] ) );
  dp_1 \layer1_reg[12][14]  ( .ip(N917), .ck(clk), .q(\layer1[12][14] ) );
  dp_1 \layer1_reg[12][13]  ( .ip(N916), .ck(clk), .q(\layer1[12][13] ) );
  dp_1 \layer1_reg[12][12]  ( .ip(N915), .ck(clk), .q(N463) );
  dp_1 \layer1_reg[11][23]  ( .ip(N911), .ck(clk), .q(\layer1[11][23] ) );
  dp_1 \layer1_reg[11][22]  ( .ip(N910), .ck(clk), .q(\layer1[11][22] ) );
  dp_1 \layer1_reg[11][21]  ( .ip(N909), .ck(clk), .q(\layer1[11][21] ) );
  dp_1 \layer1_reg[11][20]  ( .ip(N908), .ck(clk), .q(\layer1[11][20] ) );
  dp_1 \layer1_reg[11][19]  ( .ip(N907), .ck(clk), .q(\layer1[11][19] ) );
  dp_1 \layer1_reg[11][18]  ( .ip(N906), .ck(clk), .q(\layer1[11][18] ) );
  dp_1 \layer1_reg[11][17]  ( .ip(N905), .ck(clk), .q(\layer1[11][17] ) );
  dp_1 \layer1_reg[11][16]  ( .ip(N904), .ck(clk), .q(\layer1[11][16] ) );
  dp_1 \layer1_reg[11][15]  ( .ip(N903), .ck(clk), .q(\layer1[11][15] ) );
  dp_1 \layer1_reg[11][14]  ( .ip(N902), .ck(clk), .q(\layer1[11][14] ) );
  dp_1 \layer1_reg[11][13]  ( .ip(N901), .ck(clk), .q(\layer1[11][13] ) );
  dp_1 \layer1_reg[11][12]  ( .ip(N900), .ck(clk), .q(\layer1[11][12] ) );
  dp_1 \layer1_reg[11][11]  ( .ip(N899), .ck(clk), .q(\layer1[11][11] ) );
  dp_1 \layer1_reg[10][23]  ( .ip(N896), .ck(clk), .q(\layer1[10][23] ) );
  dp_1 \layer1_reg[10][22]  ( .ip(N895), .ck(clk), .q(\layer1[10][22] ) );
  dp_1 \layer1_reg[10][21]  ( .ip(N894), .ck(clk), .q(\layer1[10][21] ) );
  dp_1 \layer1_reg[10][20]  ( .ip(N893), .ck(clk), .q(\layer1[10][20] ) );
  dp_1 \layer1_reg[10][19]  ( .ip(N892), .ck(clk), .q(\layer1[10][19] ) );
  dp_1 \layer1_reg[10][18]  ( .ip(N891), .ck(clk), .q(\layer1[10][18] ) );
  dp_1 \layer1_reg[10][17]  ( .ip(N890), .ck(clk), .q(\layer1[10][17] ) );
  dp_1 \layer1_reg[10][16]  ( .ip(N889), .ck(clk), .q(\layer1[10][16] ) );
  dp_1 \layer1_reg[10][15]  ( .ip(N888), .ck(clk), .q(\layer1[10][15] ) );
  dp_1 \layer1_reg[10][14]  ( .ip(N887), .ck(clk), .q(\layer1[10][14] ) );
  dp_1 \layer1_reg[10][13]  ( .ip(N886), .ck(clk), .q(\layer1[10][13] ) );
  dp_1 \layer1_reg[10][12]  ( .ip(N885), .ck(clk), .q(\layer1[10][12] ) );
  dp_1 \layer1_reg[10][11]  ( .ip(N884), .ck(clk), .q(\layer1[10][11] ) );
  dp_1 \layer1_reg[10][10]  ( .ip(N883), .ck(clk), .q(N429) );
  dp_1 \layer1_reg[9][23]  ( .ip(N881), .ck(clk), .q(\layer1[9][23] ) );
  dp_1 \layer1_reg[9][22]  ( .ip(N880), .ck(clk), .q(\layer1[9][22] ) );
  dp_1 \layer1_reg[9][21]  ( .ip(N879), .ck(clk), .q(\layer1[9][21] ) );
  dp_1 \layer1_reg[9][20]  ( .ip(N878), .ck(clk), .q(\layer1[9][20] ) );
  dp_1 \layer1_reg[9][19]  ( .ip(N877), .ck(clk), .q(\layer1[9][19] ) );
  dp_1 \layer1_reg[9][18]  ( .ip(N876), .ck(clk), .q(\layer1[9][18] ) );
  dp_1 \layer1_reg[9][17]  ( .ip(N875), .ck(clk), .q(\layer1[9][17] ) );
  dp_1 \layer1_reg[9][16]  ( .ip(N874), .ck(clk), .q(\layer1[9][16] ) );
  dp_1 \layer1_reg[9][15]  ( .ip(N873), .ck(clk), .q(\layer1[9][15] ) );
  dp_1 \layer1_reg[9][14]  ( .ip(N872), .ck(clk), .q(\layer1[9][14] ) );
  dp_1 \layer1_reg[9][13]  ( .ip(N871), .ck(clk), .q(\layer1[9][13] ) );
  dp_1 \layer1_reg[9][12]  ( .ip(N870), .ck(clk), .q(\layer1[9][12] ) );
  dp_1 \layer1_reg[9][11]  ( .ip(N869), .ck(clk), .q(\layer1[9][11] ) );
  dp_1 \layer1_reg[9][10]  ( .ip(N868), .ck(clk), .q(\layer1[9][10] ) );
  dp_1 \layer1_reg[9][9]  ( .ip(N867), .ck(clk), .q(\layer1[9][9] ) );
  dp_1 \layer1_reg[8][23]  ( .ip(N866), .ck(clk), .q(\layer1[8][23] ) );
  dp_1 \layer1_reg[8][22]  ( .ip(N865), .ck(clk), .q(\layer1[8][22] ) );
  dp_1 \layer1_reg[8][21]  ( .ip(N864), .ck(clk), .q(\layer1[8][21] ) );
  dp_1 \layer1_reg[8][20]  ( .ip(N863), .ck(clk), .q(\layer1[8][20] ) );
  dp_1 \layer1_reg[8][19]  ( .ip(N862), .ck(clk), .q(\layer1[8][19] ) );
  dp_1 \layer1_reg[8][18]  ( .ip(N861), .ck(clk), .q(\layer1[8][18] ) );
  dp_1 \layer1_reg[8][17]  ( .ip(N860), .ck(clk), .q(\layer1[8][17] ) );
  dp_1 \layer1_reg[8][16]  ( .ip(N859), .ck(clk), .q(\layer1[8][16] ) );
  dp_1 \layer1_reg[8][15]  ( .ip(N858), .ck(clk), .q(\layer1[8][15] ) );
  dp_1 \layer1_reg[8][14]  ( .ip(N857), .ck(clk), .q(\layer1[8][14] ) );
  dp_1 \layer1_reg[8][13]  ( .ip(N856), .ck(clk), .q(\layer1[8][13] ) );
  dp_1 \layer1_reg[8][12]  ( .ip(N855), .ck(clk), .q(\layer1[8][12] ) );
  dp_1 \layer1_reg[8][11]  ( .ip(N854), .ck(clk), .q(\layer1[8][11] ) );
  dp_1 \layer1_reg[8][10]  ( .ip(N853), .ck(clk), .q(\layer1[8][10] ) );
  dp_1 \layer1_reg[8][9]  ( .ip(N852), .ck(clk), .q(\layer1[8][9] ) );
  dp_1 \layer1_reg[8][8]  ( .ip(N851), .ck(clk), .q(N395) );
  dp_1 \layer1_reg[7][22]  ( .ip(N850), .ck(clk), .q(\layer1[7][22] ) );
  dp_1 \layer1_reg[7][21]  ( .ip(N849), .ck(clk), .q(\layer1[7][21] ) );
  dp_1 \layer1_reg[7][20]  ( .ip(N848), .ck(clk), .q(\layer1[7][20] ) );
  dp_1 \layer1_reg[7][19]  ( .ip(N847), .ck(clk), .q(\layer1[7][19] ) );
  dp_1 \layer1_reg[7][18]  ( .ip(N846), .ck(clk), .q(\layer1[7][18] ) );
  dp_1 \layer1_reg[7][17]  ( .ip(N845), .ck(clk), .q(\layer1[7][17] ) );
  dp_1 \layer1_reg[7][16]  ( .ip(N844), .ck(clk), .q(\layer1[7][16] ) );
  dp_1 \layer1_reg[7][15]  ( .ip(N843), .ck(clk), .q(\layer1[7][15] ) );
  dp_1 \layer1_reg[7][14]  ( .ip(N842), .ck(clk), .q(\layer1[7][14] ) );
  dp_1 \layer1_reg[7][13]  ( .ip(N841), .ck(clk), .q(\layer1[7][13] ) );
  dp_1 \layer1_reg[7][12]  ( .ip(N840), .ck(clk), .q(\layer1[7][12] ) );
  dp_1 \layer1_reg[7][11]  ( .ip(N839), .ck(clk), .q(\layer1[7][11] ) );
  dp_1 \layer1_reg[7][10]  ( .ip(N838), .ck(clk), .q(\layer1[7][10] ) );
  dp_1 \layer1_reg[7][9]  ( .ip(N837), .ck(clk), .q(\layer1[7][9] ) );
  dp_1 \layer1_reg[7][8]  ( .ip(N836), .ck(clk), .q(\layer1[7][8] ) );
  dp_1 \layer1_reg[7][7]  ( .ip(N835), .ck(clk), .q(\layer1[7][7] ) );
  dp_1 \layer1_reg[6][21]  ( .ip(N834), .ck(clk), .q(\layer1[6][21] ) );
  dp_1 \layer1_reg[6][20]  ( .ip(N833), .ck(clk), .q(\layer1[6][20] ) );
  dp_1 \layer1_reg[6][19]  ( .ip(N832), .ck(clk), .q(\layer1[6][19] ) );
  dp_1 \layer1_reg[6][18]  ( .ip(N831), .ck(clk), .q(\layer1[6][18] ) );
  dp_1 \layer1_reg[6][17]  ( .ip(N830), .ck(clk), .q(\layer1[6][17] ) );
  dp_1 \layer1_reg[6][16]  ( .ip(N829), .ck(clk), .q(\layer1[6][16] ) );
  dp_1 \layer1_reg[6][15]  ( .ip(N828), .ck(clk), .q(\layer1[6][15] ) );
  dp_1 \layer1_reg[6][14]  ( .ip(N827), .ck(clk), .q(\layer1[6][14] ) );
  dp_1 \layer1_reg[6][13]  ( .ip(N826), .ck(clk), .q(\layer1[6][13] ) );
  dp_1 \layer1_reg[6][12]  ( .ip(N825), .ck(clk), .q(\layer1[6][12] ) );
  dp_1 \layer1_reg[6][11]  ( .ip(N824), .ck(clk), .q(\layer1[6][11] ) );
  dp_1 \layer1_reg[6][10]  ( .ip(N823), .ck(clk), .q(\layer1[6][10] ) );
  dp_1 \layer1_reg[6][9]  ( .ip(N822), .ck(clk), .q(\layer1[6][9] ) );
  dp_1 \layer1_reg[6][8]  ( .ip(N821), .ck(clk), .q(\layer1[6][8] ) );
  dp_1 \layer1_reg[6][7]  ( .ip(N820), .ck(clk), .q(\layer1[6][7] ) );
  dp_1 \layer1_reg[6][6]  ( .ip(N819), .ck(clk), .q(N361) );
  dp_1 \layer1_reg[5][20]  ( .ip(N818), .ck(clk), .q(\layer1[5][20] ) );
  dp_1 \layer1_reg[5][19]  ( .ip(N817), .ck(clk), .q(\layer1[5][19] ) );
  dp_1 \layer1_reg[5][18]  ( .ip(N816), .ck(clk), .q(\layer1[5][18] ) );
  dp_1 \layer1_reg[5][17]  ( .ip(N815), .ck(clk), .q(\layer1[5][17] ) );
  dp_1 \layer1_reg[5][16]  ( .ip(N814), .ck(clk), .q(\layer1[5][16] ) );
  dp_1 \layer1_reg[5][15]  ( .ip(N813), .ck(clk), .q(\layer1[5][15] ) );
  dp_1 \layer1_reg[5][14]  ( .ip(N812), .ck(clk), .q(\layer1[5][14] ) );
  dp_1 \layer1_reg[5][13]  ( .ip(N811), .ck(clk), .q(\layer1[5][13] ) );
  dp_1 \layer1_reg[5][12]  ( .ip(N810), .ck(clk), .q(\layer1[5][12] ) );
  dp_1 \layer1_reg[5][11]  ( .ip(N809), .ck(clk), .q(\layer1[5][11] ) );
  dp_1 \layer1_reg[5][10]  ( .ip(N808), .ck(clk), .q(\layer1[5][10] ) );
  dp_1 \layer1_reg[5][9]  ( .ip(N807), .ck(clk), .q(\layer1[5][9] ) );
  dp_1 \layer1_reg[5][8]  ( .ip(N806), .ck(clk), .q(\layer1[5][8] ) );
  dp_1 \layer1_reg[5][7]  ( .ip(N805), .ck(clk), .q(\layer1[5][7] ) );
  dp_1 \layer1_reg[5][6]  ( .ip(N804), .ck(clk), .q(\layer1[5][6] ) );
  dp_1 \layer1_reg[5][5]  ( .ip(N803), .ck(clk), .q(\layer1[5][5] ) );
  dp_1 \layer1_reg[4][19]  ( .ip(N802), .ck(clk), .q(\layer1[4][19] ) );
  dp_1 \layer1_reg[4][18]  ( .ip(N801), .ck(clk), .q(\layer1[4][18] ) );
  dp_1 \layer1_reg[4][17]  ( .ip(N800), .ck(clk), .q(\layer1[4][17] ) );
  dp_1 \layer1_reg[4][16]  ( .ip(N799), .ck(clk), .q(\layer1[4][16] ) );
  dp_1 \layer1_reg[4][15]  ( .ip(N798), .ck(clk), .q(\layer1[4][15] ) );
  dp_1 \layer1_reg[4][14]  ( .ip(N797), .ck(clk), .q(\layer1[4][14] ) );
  dp_1 \layer1_reg[4][13]  ( .ip(N796), .ck(clk), .q(\layer1[4][13] ) );
  dp_1 \layer1_reg[4][12]  ( .ip(N795), .ck(clk), .q(\layer1[4][12] ) );
  dp_1 \layer1_reg[4][11]  ( .ip(N794), .ck(clk), .q(\layer1[4][11] ) );
  dp_1 \layer1_reg[4][10]  ( .ip(N793), .ck(clk), .q(\layer1[4][10] ) );
  dp_1 \layer1_reg[4][9]  ( .ip(N792), .ck(clk), .q(\layer1[4][9] ) );
  dp_1 \layer1_reg[4][8]  ( .ip(N791), .ck(clk), .q(\layer1[4][8] ) );
  dp_1 \layer1_reg[4][7]  ( .ip(N790), .ck(clk), .q(\layer1[4][7] ) );
  dp_1 \layer1_reg[4][6]  ( .ip(N789), .ck(clk), .q(\layer1[4][6] ) );
  dp_1 \layer1_reg[4][5]  ( .ip(N788), .ck(clk), .q(\layer1[4][5] ) );
  dp_1 \layer1_reg[4][4]  ( .ip(N787), .ck(clk), .q(N327) );
  dp_1 \layer1_reg[3][18]  ( .ip(N786), .ck(clk), .q(\layer1[3][18] ) );
  dp_1 \layer1_reg[3][17]  ( .ip(N785), .ck(clk), .q(\layer1[3][17] ) );
  dp_1 \layer1_reg[3][16]  ( .ip(N784), .ck(clk), .q(\layer1[3][16] ) );
  dp_1 \layer1_reg[3][15]  ( .ip(N783), .ck(clk), .q(\layer1[3][15] ) );
  dp_1 \layer1_reg[3][14]  ( .ip(N782), .ck(clk), .q(\layer1[3][14] ) );
  dp_1 \layer1_reg[3][13]  ( .ip(N781), .ck(clk), .q(\layer1[3][13] ) );
  dp_1 \layer1_reg[3][12]  ( .ip(N780), .ck(clk), .q(\layer1[3][12] ) );
  dp_1 \layer1_reg[3][11]  ( .ip(N779), .ck(clk), .q(\layer1[3][11] ) );
  dp_1 \layer1_reg[3][10]  ( .ip(N778), .ck(clk), .q(\layer1[3][10] ) );
  dp_1 \layer1_reg[3][9]  ( .ip(N777), .ck(clk), .q(\layer1[3][9] ) );
  dp_1 \layer1_reg[3][8]  ( .ip(N776), .ck(clk), .q(\layer1[3][8] ) );
  dp_1 \layer1_reg[3][7]  ( .ip(N775), .ck(clk), .q(\layer1[3][7] ) );
  dp_1 \layer1_reg[3][6]  ( .ip(N774), .ck(clk), .q(\layer1[3][6] ) );
  dp_1 \layer1_reg[3][5]  ( .ip(N773), .ck(clk), .q(\layer1[3][5] ) );
  dp_1 \layer1_reg[3][4]  ( .ip(N772), .ck(clk), .q(\layer1[3][4] ) );
  dp_1 \layer1_reg[3][3]  ( .ip(N771), .ck(clk), .q(\layer1[3][3] ) );
  dp_1 \layer1_reg[2][17]  ( .ip(N770), .ck(clk), .q(\layer1[2][17] ) );
  dp_1 \layer1_reg[2][16]  ( .ip(N769), .ck(clk), .q(\layer1[2][16] ) );
  dp_1 \layer1_reg[2][15]  ( .ip(N768), .ck(clk), .q(\layer1[2][15] ) );
  dp_1 \layer1_reg[2][14]  ( .ip(N767), .ck(clk), .q(\layer1[2][14] ) );
  dp_1 \layer1_reg[2][13]  ( .ip(N766), .ck(clk), .q(\layer1[2][13] ) );
  dp_1 \layer1_reg[2][12]  ( .ip(N765), .ck(clk), .q(\layer1[2][12] ) );
  dp_1 \layer1_reg[2][11]  ( .ip(N764), .ck(clk), .q(\layer1[2][11] ) );
  dp_1 \layer1_reg[2][10]  ( .ip(N763), .ck(clk), .q(\layer1[2][10] ) );
  dp_1 \layer1_reg[2][9]  ( .ip(N762), .ck(clk), .q(\layer1[2][9] ) );
  dp_1 \layer1_reg[2][8]  ( .ip(N761), .ck(clk), .q(\layer1[2][8] ) );
  dp_1 \layer1_reg[2][7]  ( .ip(N760), .ck(clk), .q(\layer1[2][7] ) );
  dp_1 \layer1_reg[2][6]  ( .ip(N759), .ck(clk), .q(\layer1[2][6] ) );
  dp_1 \layer1_reg[2][5]  ( .ip(N758), .ck(clk), .q(\layer1[2][5] ) );
  dp_1 \layer1_reg[2][4]  ( .ip(N757), .ck(clk), .q(\layer1[2][4] ) );
  dp_1 \layer1_reg[2][3]  ( .ip(N756), .ck(clk), .q(\layer1[2][3] ) );
  dp_1 \layer1_reg[2][2]  ( .ip(N755), .ck(clk), .q(N293) );
  dp_1 \layer1_reg[1][16]  ( .ip(N754), .ck(clk), .q(\layer1[1][16] ) );
  dp_1 \layer1_reg[1][15]  ( .ip(N753), .ck(clk), .q(\layer1[1][15] ) );
  dp_1 \layer1_reg[1][14]  ( .ip(N752), .ck(clk), .q(\layer1[1][14] ) );
  dp_1 \layer1_reg[1][13]  ( .ip(N751), .ck(clk), .q(\layer1[1][13] ) );
  dp_1 \layer1_reg[1][12]  ( .ip(N750), .ck(clk), .q(\layer1[1][12] ) );
  dp_1 \layer1_reg[1][11]  ( .ip(N749), .ck(clk), .q(\layer1[1][11] ) );
  dp_1 \layer1_reg[1][10]  ( .ip(N748), .ck(clk), .q(\layer1[1][10] ) );
  dp_1 \layer1_reg[1][9]  ( .ip(N747), .ck(clk), .q(\layer1[1][9] ) );
  dp_1 \layer1_reg[1][8]  ( .ip(N746), .ck(clk), .q(\layer1[1][8] ) );
  dp_1 \layer1_reg[1][7]  ( .ip(N745), .ck(clk), .q(\layer1[1][7] ) );
  dp_1 \layer1_reg[1][6]  ( .ip(N744), .ck(clk), .q(\layer1[1][6] ) );
  dp_1 \layer1_reg[1][5]  ( .ip(N743), .ck(clk), .q(\layer1[1][5] ) );
  dp_1 \layer1_reg[1][4]  ( .ip(N742), .ck(clk), .q(\layer1[1][4] ) );
  dp_1 \layer1_reg[1][3]  ( .ip(N741), .ck(clk), .q(\layer1[1][3] ) );
  dp_1 \layer1_reg[1][2]  ( .ip(N740), .ck(clk), .q(\layer1[1][2] ) );
  dp_1 \layer1_reg[1][1]  ( .ip(N739), .ck(clk), .q(\layer1[1][1] ) );
  dp_1 \layer1_reg[0][16]  ( .ip(n540), .ck(clk), .q(\layer1[0][16] ) );
  dp_1 \layer1_reg[0][15]  ( .ip(N738), .ck(clk), .q(\layer1[0][15] ) );
  dp_1 \layer1_reg[0][14]  ( .ip(N737), .ck(clk), .q(\layer1[0][14] ) );
  dp_1 \layer1_reg[0][13]  ( .ip(N736), .ck(clk), .q(\layer1[0][13] ) );
  dp_1 \layer1_reg[0][12]  ( .ip(N735), .ck(clk), .q(\layer1[0][12] ) );
  dp_1 \layer1_reg[0][11]  ( .ip(N734), .ck(clk), .q(\layer1[0][11] ) );
  dp_1 \layer1_reg[0][10]  ( .ip(N733), .ck(clk), .q(\layer1[0][10] ) );
  dp_1 \layer1_reg[0][9]  ( .ip(N732), .ck(clk), .q(\layer1[0][9] ) );
  dp_1 \layer1_reg[0][8]  ( .ip(N731), .ck(clk), .q(\layer1[0][8] ) );
  dp_1 \layer1_reg[0][7]  ( .ip(N730), .ck(clk), .q(\layer1[0][7] ) );
  dp_1 \layer1_reg[0][6]  ( .ip(N729), .ck(clk), .q(\layer1[0][6] ) );
  dp_1 \layer1_reg[0][5]  ( .ip(N728), .ck(clk), .q(\layer1[0][5] ) );
  dp_1 \layer1_reg[0][4]  ( .ip(N727), .ck(clk), .q(\layer1[0][4] ) );
  dp_1 \layer1_reg[0][3]  ( .ip(N726), .ck(clk), .q(\layer1[0][3] ) );
  dp_1 \layer1_reg[0][2]  ( .ip(N725), .ck(clk), .q(\layer1[0][2] ) );
  dp_1 \layer1_reg[0][1]  ( .ip(N724), .ck(clk), .q(\layer1[0][1] ) );
  buf_1 U765 ( .ip(reset), .op(n483) );
  or2_1 U766 ( .ip1(w[15]), .ip2(n483), .op(n293) );
  or2_1 U767 ( .ip1(in[8]), .ip2(n483), .op(n284) );
  nand2_1 U768 ( .ip1(n293), .ip2(n284), .op(N971) );
  or2_1 U769 ( .ip1(in[7]), .ip2(n483), .op(n285) );
  nand2_1 U770 ( .ip1(n293), .ip2(n285), .op(N970) );
  or2_1 U771 ( .ip1(in[6]), .ip2(n483), .op(n286) );
  nand2_1 U772 ( .ip1(n293), .ip2(n286), .op(N969) );
  or2_1 U773 ( .ip1(in[5]), .ip2(n483), .op(n287) );
  nand2_1 U774 ( .ip1(n293), .ip2(n287), .op(N968) );
  or2_1 U775 ( .ip1(in[4]), .ip2(n483), .op(n288) );
  nand2_1 U776 ( .ip1(n293), .ip2(n288), .op(N967) );
  or2_1 U777 ( .ip1(in[3]), .ip2(n483), .op(n289) );
  nand2_1 U778 ( .ip1(n293), .ip2(n289), .op(N966) );
  or2_1 U779 ( .ip1(in[2]), .ip2(n483), .op(n290) );
  nand2_1 U780 ( .ip1(n293), .ip2(n290), .op(N965) );
  or2_1 U781 ( .ip1(in[1]), .ip2(reset), .op(n291) );
  nand2_1 U782 ( .ip1(n293), .ip2(n291), .op(N964) );
  or2_1 U783 ( .ip1(in[0]), .ip2(n483), .op(n292) );
  nand2_1 U784 ( .ip1(n293), .ip2(n292), .op(N963) );
  or2_1 U785 ( .ip1(in[15]), .ip2(n483), .op(n303) );
  or2_1 U786 ( .ip1(w[8]), .ip2(n483), .op(n294) );
  nand2_1 U787 ( .ip1(n303), .ip2(n294), .op(N866) );
  or2_1 U788 ( .ip1(w[7]), .ip2(n483), .op(n295) );
  nand2_1 U789 ( .ip1(n303), .ip2(n295), .op(N850) );
  or2_1 U790 ( .ip1(w[6]), .ip2(reset), .op(n296) );
  nand2_1 U791 ( .ip1(n303), .ip2(n296), .op(N834) );
  or2_1 U792 ( .ip1(w[5]), .ip2(reset), .op(n297) );
  nand2_1 U793 ( .ip1(n303), .ip2(n297), .op(N818) );
  or2_1 U794 ( .ip1(w[4]), .ip2(n483), .op(n298) );
  nand2_1 U795 ( .ip1(n303), .ip2(n298), .op(N802) );
  or2_1 U796 ( .ip1(w[3]), .ip2(reset), .op(n299) );
  nand2_1 U797 ( .ip1(n303), .ip2(n299), .op(N786) );
  or2_1 U798 ( .ip1(w[2]), .ip2(reset), .op(n300) );
  nand2_1 U799 ( .ip1(n303), .ip2(n300), .op(N770) );
  or2_1 U800 ( .ip1(w[1]), .ip2(reset), .op(n301) );
  nand2_1 U801 ( .ip1(n303), .ip2(n301), .op(N754) );
  or2_1 U802 ( .ip1(w[0]), .ip2(n483), .op(n302) );
  nand2_1 U803 ( .ip1(n303), .ip2(n302), .op(N738) );
  nand2_1 U804 ( .ip1(\layer3[1][5] ), .ip2(\layer3[0][5] ), .op(n306) );
  or2_1 U805 ( .ip1(\layer3[1][5] ), .ip2(\layer3[0][5] ), .op(n304) );
  nand3_1 U806 ( .ip1(\layer3[1][4] ), .ip2(\layer3[0][4] ), .ip3(n304), .op(
        n305) );
  nand2_1 U807 ( .ip1(n306), .ip2(n305), .op(n307) );
  fulladder U808 ( .a(\layer3[1][6] ), .b(\layer3[0][6] ), .ci(n307), .co(n308), .s() );
  fulladder U809 ( .a(\layer3[1][7] ), .b(\layer3[0][7] ), .ci(n308), .co(n310), .s() );
  inv_1 U810 ( .ip(reset), .op(n778) );
  and2_1 U811 ( .ip1(n309), .ip2(n778), .op(N1371) );
  fulladder U812 ( .a(\layer3[1][8] ), .b(\layer3[0][8] ), .ci(n310), .co(n312), .s(n309) );
  and2_1 U813 ( .ip1(n311), .ip2(n778), .op(N1372) );
  fulladder U814 ( .a(\layer3[1][9] ), .b(\layer3[0][9] ), .ci(n312), .co(n314), .s(n311) );
  inv_1 U815 ( .ip(reset), .op(n835) );
  and2_1 U816 ( .ip1(n313), .ip2(n835), .op(N1373) );
  fulladder U817 ( .a(\layer3[1][10] ), .b(\layer3[0][10] ), .ci(n314), .co(
        n316), .s(n313) );
  and2_1 U818 ( .ip1(n315), .ip2(n835), .op(N1374) );
  fulladder U819 ( .a(\layer3[1][11] ), .b(\layer3[0][11] ), .ci(n316), .co(
        n318), .s(n315) );
  and2_1 U820 ( .ip1(n317), .ip2(n835), .op(N1375) );
  fulladder U821 ( .a(\layer3[1][12] ), .b(\layer3[0][12] ), .ci(n318), .co(
        n320), .s(n317) );
  and2_1 U822 ( .ip1(n319), .ip2(n835), .op(N1376) );
  fulladder U823 ( .a(\layer3[1][13] ), .b(\layer3[0][13] ), .ci(n320), .co(
        n322), .s(n319) );
  and2_1 U824 ( .ip1(n321), .ip2(n835), .op(N1377) );
  fulladder U825 ( .a(\layer3[1][14] ), .b(\layer3[0][14] ), .ci(n322), .co(
        n324), .s(n321) );
  and2_1 U826 ( .ip1(n323), .ip2(n835), .op(N1378) );
  fulladder U827 ( .a(\layer3[1][15] ), .b(\layer3[0][15] ), .ci(n324), .co(
        n326), .s(n323) );
  and2_1 U828 ( .ip1(n325), .ip2(n835), .op(N1379) );
  fulladder U829 ( .a(\layer3[1][16] ), .b(\layer3[0][16] ), .ci(n326), .co(
        n328), .s(n325) );
  and2_1 U830 ( .ip1(n327), .ip2(n835), .op(N1380) );
  fulladder U831 ( .a(\layer3[1][17] ), .b(\layer3[0][17] ), .ci(n328), .co(
        n330), .s(n327) );
  and2_1 U832 ( .ip1(n329), .ip2(n835), .op(N1381) );
  fulladder U833 ( .a(\layer3[1][18] ), .b(\layer3[0][18] ), .ci(n330), .co(
        n332), .s(n329) );
  and2_1 U834 ( .ip1(n331), .ip2(n835), .op(N1382) );
  fulladder U835 ( .a(\layer3[1][19] ), .b(\layer3[0][19] ), .ci(n332), .co(
        n334), .s(n331) );
  and2_1 U836 ( .ip1(n333), .ip2(n835), .op(N1383) );
  fulladder U837 ( .a(\layer3[1][20] ), .b(\layer3[0][20] ), .ci(n334), .co(
        n337), .s(n333) );
  nor2_1 U838 ( .ip1(n337), .ip2(\layer3[1][21] ), .op(n336) );
  nand2_1 U839 ( .ip1(n337), .ip2(\layer3[1][21] ), .op(n339) );
  inv_1 U840 ( .ip(n339), .op(n335) );
  nor3_1 U841 ( .ip1(n336), .ip2(n483), .ip3(n335), .op(N1384) );
  inv_1 U842 ( .ip(\layer3[1][22] ), .op(n338) );
  and3_1 U843 ( .ip1(n337), .ip2(\layer3[1][21] ), .ip3(\layer3[1][22] ), .op(
        n341) );
  not_ab_or_c_or_d U844 ( .ip1(n339), .ip2(n338), .ip3(reset), .ip4(n341), 
        .op(N1385) );
  nor2_1 U845 ( .ip1(\layer3[1][23] ), .ip2(n341), .op(n340) );
  not_ab_or_c_or_d U846 ( .ip1(\layer3[1][23] ), .ip2(n341), .ip3(reset), 
        .ip4(n340), .op(N1386) );
  and2_1 U847 ( .ip1(N675), .ip2(n835), .op(N1395) );
  and2_1 U848 ( .ip1(N676), .ip2(n801), .op(N1396) );
  and2_1 U849 ( .ip1(N677), .ip2(n778), .op(N1397) );
  and2_1 U850 ( .ip1(N678), .ip2(n672), .op(N1398) );
  nor2_1 U851 ( .ip1(\layer3[2][12] ), .ip2(\layer3[3][12] ), .op(n342) );
  nand2_1 U852 ( .ip1(\layer3[2][12] ), .ip2(\layer3[3][12] ), .op(n343) );
  inv_1 U853 ( .ip(n343), .op(n344) );
  nor3_1 U854 ( .ip1(n342), .ip2(n483), .ip3(n344), .op(N1399) );
  mux2_1 U855 ( .ip1(n344), .ip2(n343), .s(\layer3[3][13] ), .op(n346) );
  nor2_1 U856 ( .ip1(\layer3[2][13] ), .ip2(n346), .op(n345) );
  not_ab_or_c_or_d U857 ( .ip1(\layer3[2][13] ), .ip2(n346), .ip3(reset), 
        .ip4(n345), .op(N1400) );
  nand2_1 U858 ( .ip1(\layer3[3][13] ), .ip2(\layer3[2][13] ), .op(n349) );
  or2_1 U859 ( .ip1(\layer3[3][13] ), .ip2(\layer3[2][13] ), .op(n347) );
  nand3_1 U860 ( .ip1(\layer3[3][12] ), .ip2(\layer3[2][12] ), .ip3(n347), 
        .op(n348) );
  nand2_1 U861 ( .ip1(n349), .ip2(n348), .op(n351) );
  and2_1 U862 ( .ip1(n350), .ip2(n778), .op(N1401) );
  fulladder U863 ( .a(\layer3[3][14] ), .b(\layer3[2][14] ), .ci(n351), .co(
        n353), .s(n350) );
  and2_1 U864 ( .ip1(n352), .ip2(n801), .op(N1402) );
  fulladder U865 ( .a(\layer3[3][15] ), .b(\layer3[2][15] ), .ci(n353), .co(
        n355), .s(n352) );
  and2_1 U866 ( .ip1(n354), .ip2(n778), .op(N1403) );
  fulladder U867 ( .a(\layer3[3][16] ), .b(\layer3[2][16] ), .ci(n355), .co(
        n357), .s(n354) );
  and2_1 U868 ( .ip1(n356), .ip2(n801), .op(N1404) );
  fulladder U869 ( .a(\layer3[3][17] ), .b(\layer3[2][17] ), .ci(n357), .co(
        n359), .s(n356) );
  and2_1 U870 ( .ip1(n358), .ip2(n778), .op(N1405) );
  fulladder U871 ( .a(\layer3[3][18] ), .b(\layer3[2][18] ), .ci(n359), .co(
        n361), .s(n358) );
  and2_1 U872 ( .ip1(n360), .ip2(n835), .op(N1406) );
  fulladder U873 ( .a(\layer3[3][19] ), .b(\layer3[2][19] ), .ci(n361), .co(
        n363), .s(n360) );
  and2_1 U874 ( .ip1(n362), .ip2(n672), .op(N1407) );
  fulladder U875 ( .a(\layer3[3][20] ), .b(\layer3[2][20] ), .ci(n363), .co(
        n365), .s(n362) );
  and2_1 U876 ( .ip1(n364), .ip2(n672), .op(N1408) );
  fulladder U877 ( .a(\layer3[3][21] ), .b(\layer3[2][21] ), .ci(n365), .co(
        n367), .s(n364) );
  and2_1 U878 ( .ip1(n366), .ip2(n672), .op(N1409) );
  fulladder U879 ( .a(\layer3[3][22] ), .b(\layer3[2][22] ), .ci(n367), .co(
        n370), .s(n366) );
  xor2_1 U880 ( .ip1(\layer3[3][23] ), .ip2(\layer3[2][23] ), .op(n369) );
  nor2_1 U881 ( .ip1(n370), .ip2(n369), .op(n368) );
  not_ab_or_c_or_d U882 ( .ip1(n370), .ip2(n369), .ip3(reset), .ip4(n368), 
        .op(N1410) );
  nand2_1 U883 ( .ip1(\layer2[1][3] ), .ip2(\layer2[0][3] ), .op(n373) );
  or2_1 U884 ( .ip1(\layer2[1][3] ), .ip2(\layer2[0][3] ), .op(n371) );
  nand3_1 U885 ( .ip1(\layer2[1][2] ), .ip2(\layer2[0][2] ), .ip3(n371), .op(
        n372) );
  nand2_1 U886 ( .ip1(n373), .ip2(n372), .op(n375) );
  inv_1 U887 ( .ip(reset), .op(n540) );
  and2_1 U888 ( .ip1(n374), .ip2(n540), .op(N1239) );
  fulladder U889 ( .a(\layer2[1][4] ), .b(\layer2[0][4] ), .ci(n375), .co(n377), .s(n374) );
  and2_1 U890 ( .ip1(n376), .ip2(n540), .op(N1240) );
  fulladder U891 ( .a(\layer2[1][5] ), .b(\layer2[0][5] ), .ci(n377), .co(n379), .s(n376) );
  and2_1 U892 ( .ip1(n378), .ip2(n540), .op(N1241) );
  fulladder U893 ( .a(\layer2[1][6] ), .b(\layer2[0][6] ), .ci(n379), .co(n381), .s(n378) );
  and2_1 U894 ( .ip1(n380), .ip2(n540), .op(N1242) );
  fulladder U895 ( .a(\layer2[1][7] ), .b(\layer2[0][7] ), .ci(n381), .co(n383), .s(n380) );
  and2_1 U896 ( .ip1(n382), .ip2(n540), .op(N1243) );
  fulladder U897 ( .a(\layer2[1][8] ), .b(\layer2[0][8] ), .ci(n383), .co(n385), .s(n382) );
  and2_1 U898 ( .ip1(n384), .ip2(n540), .op(N1244) );
  fulladder U899 ( .a(\layer2[1][9] ), .b(\layer2[0][9] ), .ci(n385), .co(n387), .s(n384) );
  and2_1 U900 ( .ip1(n386), .ip2(n540), .op(N1245) );
  fulladder U901 ( .a(\layer2[1][10] ), .b(\layer2[0][10] ), .ci(n387), .co(
        n389), .s(n386) );
  and2_1 U902 ( .ip1(n388), .ip2(n540), .op(N1246) );
  fulladder U903 ( .a(\layer2[1][11] ), .b(\layer2[0][11] ), .ci(n389), .co(
        n391), .s(n388) );
  and2_1 U904 ( .ip1(n390), .ip2(n540), .op(N1247) );
  fulladder U905 ( .a(\layer2[1][12] ), .b(\layer2[0][12] ), .ci(n391), .co(
        n393), .s(n390) );
  and2_1 U906 ( .ip1(n392), .ip2(n540), .op(N1248) );
  fulladder U907 ( .a(\layer2[1][13] ), .b(\layer2[0][13] ), .ci(n393), .co(
        n395), .s(n392) );
  and2_1 U908 ( .ip1(n394), .ip2(n540), .op(N1249) );
  fulladder U909 ( .a(\layer2[1][14] ), .b(\layer2[0][14] ), .ci(n395), .co(
        n397), .s(n394) );
  and2_1 U910 ( .ip1(n396), .ip2(n540), .op(N1250) );
  fulladder U911 ( .a(\layer2[1][15] ), .b(\layer2[0][15] ), .ci(n397), .co(
        n399), .s(n396) );
  and2_1 U912 ( .ip1(n398), .ip2(n540), .op(N1251) );
  fulladder U913 ( .a(\layer2[1][16] ), .b(\layer2[0][16] ), .ci(n399), .co(
        n401), .s(n398) );
  and2_1 U914 ( .ip1(n400), .ip2(n540), .op(N1252) );
  fulladder U915 ( .a(\layer2[1][17] ), .b(\layer2[0][17] ), .ci(n401), .co(
        n404), .s(n400) );
  nor2_1 U916 ( .ip1(n404), .ip2(\layer2[1][18] ), .op(n403) );
  nand2_1 U917 ( .ip1(n404), .ip2(\layer2[1][18] ), .op(n407) );
  inv_1 U918 ( .ip(n407), .op(n402) );
  nor3_1 U919 ( .ip1(n403), .ip2(n483), .ip3(n402), .op(N1253) );
  inv_1 U920 ( .ip(\layer2[1][19] ), .op(n406) );
  and3_1 U921 ( .ip1(n404), .ip2(\layer2[1][18] ), .ip3(\layer2[1][19] ), .op(
        n405) );
  not_ab_or_c_or_d U922 ( .ip1(n407), .ip2(n406), .ip3(reset), .ip4(n405), 
        .op(N1254) );
  nor3_1 U923 ( .ip1(reset), .ip2(n407), .ip3(n406), .op(N1255) );
  and2_1 U924 ( .ip1(N551), .ip2(n540), .op(N1271) );
  and2_1 U925 ( .ip1(N552), .ip2(n540), .op(N1272) );
  nor2_1 U926 ( .ip1(\layer2[2][6] ), .ip2(\layer2[3][6] ), .op(n408) );
  nand2_1 U927 ( .ip1(\layer2[2][6] ), .ip2(\layer2[3][6] ), .op(n409) );
  inv_1 U928 ( .ip(n409), .op(n410) );
  nor3_1 U929 ( .ip1(n408), .ip2(n483), .ip3(n410), .op(N1273) );
  mux2_1 U930 ( .ip1(n410), .ip2(n409), .s(\layer2[3][7] ), .op(n412) );
  nor2_1 U931 ( .ip1(\layer2[2][7] ), .ip2(n412), .op(n411) );
  not_ab_or_c_or_d U932 ( .ip1(\layer2[2][7] ), .ip2(n412), .ip3(reset), .ip4(
        n411), .op(N1274) );
  nand2_1 U933 ( .ip1(\layer2[3][7] ), .ip2(\layer2[2][7] ), .op(n415) );
  or2_1 U934 ( .ip1(\layer2[3][7] ), .ip2(\layer2[2][7] ), .op(n413) );
  nand3_1 U935 ( .ip1(\layer2[3][6] ), .ip2(\layer2[2][6] ), .ip3(n413), .op(
        n414) );
  nand2_1 U936 ( .ip1(n415), .ip2(n414), .op(n417) );
  and2_1 U937 ( .ip1(n416), .ip2(n540), .op(N1275) );
  fulladder U938 ( .a(\layer2[3][8] ), .b(\layer2[2][8] ), .ci(n417), .co(n419), .s(n416) );
  and2_1 U939 ( .ip1(n418), .ip2(n540), .op(N1276) );
  fulladder U940 ( .a(\layer2[3][9] ), .b(\layer2[2][9] ), .ci(n419), .co(n421), .s(n418) );
  and2_1 U941 ( .ip1(n420), .ip2(n540), .op(N1277) );
  fulladder U942 ( .a(\layer2[3][10] ), .b(\layer2[2][10] ), .ci(n421), .co(
        n423), .s(n420) );
  and2_1 U943 ( .ip1(n422), .ip2(n540), .op(N1278) );
  fulladder U944 ( .a(\layer2[3][11] ), .b(\layer2[2][11] ), .ci(n423), .co(
        n425), .s(n422) );
  and2_1 U945 ( .ip1(n424), .ip2(n540), .op(N1279) );
  fulladder U946 ( .a(\layer2[3][12] ), .b(\layer2[2][12] ), .ci(n425), .co(
        n427), .s(n424) );
  and2_1 U947 ( .ip1(n426), .ip2(n540), .op(N1280) );
  fulladder U948 ( .a(\layer2[3][13] ), .b(\layer2[2][13] ), .ci(n427), .co(
        n429), .s(n426) );
  and2_1 U949 ( .ip1(n428), .ip2(n540), .op(N1281) );
  fulladder U950 ( .a(\layer2[3][14] ), .b(\layer2[2][14] ), .ci(n429), .co(
        n431), .s(n428) );
  and2_1 U951 ( .ip1(n430), .ip2(n540), .op(N1282) );
  fulladder U952 ( .a(\layer2[3][15] ), .b(\layer2[2][15] ), .ci(n431), .co(
        n433), .s(n430) );
  and2_1 U953 ( .ip1(n432), .ip2(n778), .op(N1283) );
  fulladder U954 ( .a(\layer2[3][16] ), .b(\layer2[2][16] ), .ci(n433), .co(
        n435), .s(n432) );
  and2_1 U955 ( .ip1(n434), .ip2(n778), .op(N1284) );
  fulladder U956 ( .a(\layer2[3][17] ), .b(\layer2[2][17] ), .ci(n435), .co(
        n437), .s(n434) );
  and2_1 U957 ( .ip1(n436), .ip2(n778), .op(N1285) );
  fulladder U958 ( .a(\layer2[3][18] ), .b(\layer2[2][18] ), .ci(n437), .co(
        n439), .s(n436) );
  and2_1 U959 ( .ip1(n438), .ip2(n778), .op(N1286) );
  fulladder U960 ( .a(\layer2[3][19] ), .b(\layer2[2][19] ), .ci(n439), .co(
        n441), .s(n438) );
  and2_1 U961 ( .ip1(n440), .ip2(n778), .op(N1287) );
  fulladder U962 ( .a(\layer2[3][20] ), .b(\layer2[2][20] ), .ci(n441), .co(
        n443), .s(n440) );
  and2_1 U963 ( .ip1(n442), .ip2(n778), .op(N1288) );
  fulladder U964 ( .a(\layer2[3][21] ), .b(\layer2[2][21] ), .ci(n443), .co(
        n446), .s(n442) );
  nor2_1 U965 ( .ip1(n446), .ip2(\layer2[3][22] ), .op(n445) );
  nand2_1 U966 ( .ip1(n446), .ip2(\layer2[3][22] ), .op(n449) );
  inv_1 U967 ( .ip(n449), .op(n444) );
  nor3_1 U968 ( .ip1(n445), .ip2(n483), .ip3(n444), .op(N1289) );
  inv_1 U969 ( .ip(\layer2[3][23] ), .op(n448) );
  and3_1 U970 ( .ip1(n446), .ip2(\layer2[3][22] ), .ip3(\layer2[3][23] ), .op(
        n447) );
  not_ab_or_c_or_d U971 ( .ip1(n449), .ip2(n448), .ip3(reset), .ip4(n447), 
        .op(N1290) );
  and2_1 U972 ( .ip1(N587), .ip2(n778), .op(N1307) );
  and2_1 U973 ( .ip1(N588), .ip2(n778), .op(N1308) );
  nor2_1 U974 ( .ip1(\layer2[4][10] ), .ip2(\layer2[5][10] ), .op(n450) );
  nand2_1 U975 ( .ip1(\layer2[4][10] ), .ip2(\layer2[5][10] ), .op(n451) );
  inv_1 U976 ( .ip(n451), .op(n452) );
  nor3_1 U977 ( .ip1(n450), .ip2(n483), .ip3(n452), .op(N1309) );
  mux2_1 U978 ( .ip1(n452), .ip2(n451), .s(\layer2[5][11] ), .op(n454) );
  nor2_1 U979 ( .ip1(\layer2[4][11] ), .ip2(n454), .op(n453) );
  not_ab_or_c_or_d U980 ( .ip1(\layer2[4][11] ), .ip2(n454), .ip3(reset), 
        .ip4(n453), .op(N1310) );
  nand2_1 U981 ( .ip1(\layer2[5][11] ), .ip2(\layer2[4][11] ), .op(n457) );
  or2_1 U982 ( .ip1(\layer2[5][11] ), .ip2(\layer2[4][11] ), .op(n455) );
  nand3_1 U983 ( .ip1(\layer2[5][10] ), .ip2(\layer2[4][10] ), .ip3(n455), 
        .op(n456) );
  nand2_1 U984 ( .ip1(n457), .ip2(n456), .op(n459) );
  and2_1 U985 ( .ip1(n458), .ip2(n778), .op(N1311) );
  fulladder U986 ( .a(\layer2[5][12] ), .b(\layer2[4][12] ), .ci(n459), .co(
        n461), .s(n458) );
  and2_1 U987 ( .ip1(n460), .ip2(n778), .op(N1312) );
  fulladder U988 ( .a(\layer2[5][13] ), .b(\layer2[4][13] ), .ci(n461), .co(
        n463), .s(n460) );
  and2_1 U989 ( .ip1(n462), .ip2(n778), .op(N1313) );
  fulladder U990 ( .a(\layer2[5][14] ), .b(\layer2[4][14] ), .ci(n463), .co(
        n465), .s(n462) );
  inv_1 U991 ( .ip(reset), .op(n801) );
  and2_1 U992 ( .ip1(n464), .ip2(n801), .op(N1314) );
  fulladder U993 ( .a(\layer2[5][15] ), .b(\layer2[4][15] ), .ci(n465), .co(
        n467), .s(n464) );
  and2_1 U994 ( .ip1(n466), .ip2(n801), .op(N1315) );
  fulladder U995 ( .a(\layer2[5][16] ), .b(\layer2[4][16] ), .ci(n467), .co(
        n469), .s(n466) );
  and2_1 U996 ( .ip1(n468), .ip2(n801), .op(N1316) );
  fulladder U997 ( .a(\layer2[5][17] ), .b(\layer2[4][17] ), .ci(n469), .co(
        n471), .s(n468) );
  and2_1 U998 ( .ip1(n470), .ip2(n801), .op(N1317) );
  fulladder U999 ( .a(\layer2[5][18] ), .b(\layer2[4][18] ), .ci(n471), .co(
        n473), .s(n470) );
  and2_1 U1000 ( .ip1(n472), .ip2(n801), .op(N1318) );
  fulladder U1001 ( .a(\layer2[5][19] ), .b(\layer2[4][19] ), .ci(n473), .co(
        n475), .s(n472) );
  and2_1 U1002 ( .ip1(n474), .ip2(n801), .op(N1319) );
  fulladder U1003 ( .a(\layer2[5][20] ), .b(\layer2[4][20] ), .ci(n475), .co(
        n477), .s(n474) );
  and2_1 U1004 ( .ip1(n476), .ip2(n801), .op(N1320) );
  fulladder U1005 ( .a(\layer2[5][21] ), .b(\layer2[4][21] ), .ci(n477), .co(
        n479), .s(n476) );
  and2_1 U1006 ( .ip1(n478), .ip2(n801), .op(N1321) );
  fulladder U1007 ( .a(\layer2[5][22] ), .b(\layer2[4][22] ), .ci(n479), .co(
        n482), .s(n478) );
  xor2_1 U1008 ( .ip1(\layer2[4][23] ), .ip2(\layer2[5][23] ), .op(n481) );
  nor2_1 U1009 ( .ip1(n482), .ip2(n481), .op(n480) );
  not_ab_or_c_or_d U1010 ( .ip1(n482), .ip2(n481), .ip3(reset), .ip4(n480), 
        .op(N1322) );
  and2_1 U1011 ( .ip1(N623), .ip2(n801), .op(N1343) );
  and2_1 U1012 ( .ip1(N624), .ip2(n801), .op(N1344) );
  nor2_1 U1013 ( .ip1(\layer2[6][14] ), .ip2(\layer2[7][14] ), .op(n484) );
  nand2_1 U1014 ( .ip1(\layer2[6][14] ), .ip2(\layer2[7][14] ), .op(n485) );
  inv_1 U1015 ( .ip(n485), .op(n486) );
  nor3_1 U1016 ( .ip1(n484), .ip2(n483), .ip3(n486), .op(N1345) );
  mux2_1 U1017 ( .ip1(n486), .ip2(n485), .s(\layer2[7][15] ), .op(n488) );
  nor2_1 U1018 ( .ip1(\layer2[6][15] ), .ip2(n488), .op(n487) );
  not_ab_or_c_or_d U1019 ( .ip1(\layer2[6][15] ), .ip2(n488), .ip3(reset), 
        .ip4(n487), .op(N1346) );
  nand2_1 U1020 ( .ip1(\layer2[7][15] ), .ip2(\layer2[6][15] ), .op(n491) );
  or2_1 U1021 ( .ip1(\layer2[7][15] ), .ip2(\layer2[6][15] ), .op(n489) );
  nand3_1 U1022 ( .ip1(\layer2[7][14] ), .ip2(\layer2[6][14] ), .ip3(n489), 
        .op(n490) );
  nand2_1 U1023 ( .ip1(n491), .ip2(n490), .op(n493) );
  and2_1 U1024 ( .ip1(n492), .ip2(n801), .op(N1347) );
  fulladder U1025 ( .a(\layer2[7][16] ), .b(\layer2[6][16] ), .ci(n493), .co(
        n495), .s(n492) );
  and2_1 U1026 ( .ip1(n494), .ip2(n540), .op(N1348) );
  fulladder U1027 ( .a(\layer2[7][17] ), .b(\layer2[6][17] ), .ci(n495), .co(
        n497), .s(n494) );
  and2_1 U1028 ( .ip1(n496), .ip2(n801), .op(N1349) );
  fulladder U1029 ( .a(\layer2[7][18] ), .b(\layer2[6][18] ), .ci(n497), .co(
        n499), .s(n496) );
  and2_1 U1030 ( .ip1(n498), .ip2(n540), .op(N1350) );
  fulladder U1031 ( .a(\layer2[7][19] ), .b(\layer2[6][19] ), .ci(n499), .co(
        n501), .s(n498) );
  and2_1 U1032 ( .ip1(n500), .ip2(n540), .op(N1351) );
  fulladder U1033 ( .a(\layer2[7][20] ), .b(\layer2[6][20] ), .ci(n501), .co(
        n503), .s(n500) );
  and2_1 U1034 ( .ip1(n502), .ip2(n540), .op(N1352) );
  fulladder U1035 ( .a(\layer2[7][21] ), .b(\layer2[6][21] ), .ci(n503), .co(
        n505), .s(n502) );
  and2_1 U1036 ( .ip1(n504), .ip2(n540), .op(N1353) );
  fulladder U1037 ( .a(\layer2[7][22] ), .b(\layer2[6][22] ), .ci(n505), .co(
        n508), .s(n504) );
  xor2_1 U1038 ( .ip1(\layer2[6][23] ), .ip2(\layer2[7][23] ), .op(n507) );
  nor2_1 U1039 ( .ip1(n508), .ip2(n507), .op(n506) );
  not_ab_or_c_or_d U1040 ( .ip1(n508), .ip2(n507), .ip3(reset), .ip4(n506), 
        .op(N1354) );
  nand2_1 U1041 ( .ip1(\layer1[1][1] ), .ip2(\layer1[0][1] ), .op(n509) );
  inv_1 U1042 ( .ip(n509), .op(n510) );
  mux2_1 U1043 ( .ip1(n510), .ip2(n509), .s(\layer1[0][2] ), .op(n512) );
  nor2_1 U1044 ( .ip1(\layer1[1][2] ), .ip2(n512), .op(n511) );
  not_ab_or_c_or_d U1045 ( .ip1(\layer1[1][2] ), .ip2(n512), .ip3(reset), 
        .ip4(n511), .op(N981) );
  nand2_1 U1046 ( .ip1(\layer1[0][2] ), .ip2(\layer1[1][2] ), .op(n515) );
  or2_1 U1047 ( .ip1(\layer1[0][2] ), .ip2(\layer1[1][2] ), .op(n513) );
  nand3_1 U1048 ( .ip1(\layer1[0][1] ), .ip2(\layer1[1][1] ), .ip3(n513), .op(
        n514) );
  nand2_1 U1049 ( .ip1(n515), .ip2(n514), .op(n517) );
  and2_1 U1050 ( .ip1(n516), .ip2(n540), .op(N982) );
  fulladder U1051 ( .a(\layer1[0][3] ), .b(\layer1[1][3] ), .ci(n517), .co(
        n519), .s(n516) );
  and2_1 U1052 ( .ip1(n518), .ip2(n540), .op(N983) );
  fulladder U1053 ( .a(\layer1[0][4] ), .b(\layer1[1][4] ), .ci(n519), .co(
        n521), .s(n518) );
  and2_1 U1054 ( .ip1(n520), .ip2(n540), .op(N984) );
  fulladder U1055 ( .a(\layer1[0][5] ), .b(\layer1[1][5] ), .ci(n521), .co(
        n523), .s(n520) );
  and2_1 U1056 ( .ip1(n522), .ip2(n540), .op(N985) );
  fulladder U1057 ( .a(\layer1[0][6] ), .b(\layer1[1][6] ), .ci(n523), .co(
        n525), .s(n522) );
  and2_1 U1058 ( .ip1(n524), .ip2(n540), .op(N986) );
  fulladder U1059 ( .a(\layer1[0][7] ), .b(\layer1[1][7] ), .ci(n525), .co(
        n527), .s(n524) );
  and2_1 U1060 ( .ip1(n526), .ip2(n540), .op(N987) );
  fulladder U1061 ( .a(\layer1[0][8] ), .b(\layer1[1][8] ), .ci(n527), .co(
        n529), .s(n526) );
  and2_1 U1062 ( .ip1(n528), .ip2(n778), .op(N988) );
  fulladder U1063 ( .a(\layer1[0][9] ), .b(\layer1[1][9] ), .ci(n529), .co(
        n531), .s(n528) );
  and2_1 U1064 ( .ip1(n530), .ip2(n778), .op(N989) );
  fulladder U1065 ( .a(\layer1[0][10] ), .b(\layer1[1][10] ), .ci(n531), .co(
        n533), .s(n530) );
  and2_1 U1066 ( .ip1(n532), .ip2(n778), .op(N990) );
  fulladder U1067 ( .a(\layer1[0][11] ), .b(\layer1[1][11] ), .ci(n533), .co(
        n535), .s(n532) );
  and2_1 U1068 ( .ip1(n534), .ip2(n778), .op(N991) );
  fulladder U1069 ( .a(\layer1[0][12] ), .b(\layer1[1][12] ), .ci(n535), .co(
        n537), .s(n534) );
  and2_1 U1070 ( .ip1(n536), .ip2(n778), .op(N992) );
  fulladder U1071 ( .a(\layer1[0][13] ), .b(\layer1[1][13] ), .ci(n537), .co(
        n539), .s(n536) );
  and2_1 U1072 ( .ip1(n538), .ip2(n778), .op(N993) );
  fulladder U1073 ( .a(\layer1[0][14] ), .b(\layer1[1][14] ), .ci(n539), .co(
        n542), .s(n538) );
  and2_1 U1074 ( .ip1(n541), .ip2(n540), .op(N994) );
  fulladder U1075 ( .a(\layer1[0][15] ), .b(\layer1[1][15] ), .ci(n542), .co(
        n544), .s(n541) );
  and2_1 U1076 ( .ip1(n543), .ip2(n778), .op(N995) );
  fulladder U1077 ( .a(\layer1[0][16] ), .b(\layer1[1][16] ), .ci(n544), .co(
        n545), .s(n543) );
  and2_1 U1078 ( .ip1(n545), .ip2(n778), .op(N996) );
  and2_1 U1079 ( .ip1(N293), .ip2(n778), .op(N1013) );
  nor2_1 U1080 ( .ip1(\layer1[3][3] ), .ip2(\layer1[2][3] ), .op(n546) );
  nand2_1 U1081 ( .ip1(\layer1[3][3] ), .ip2(\layer1[2][3] ), .op(n547) );
  inv_1 U1082 ( .ip(n547), .op(n548) );
  nor3_1 U1083 ( .ip1(n546), .ip2(n483), .ip3(n548), .op(N1014) );
  mux2_1 U1084 ( .ip1(n548), .ip2(n547), .s(\layer1[2][4] ), .op(n550) );
  nor2_1 U1085 ( .ip1(\layer1[3][4] ), .ip2(n550), .op(n549) );
  not_ab_or_c_or_d U1086 ( .ip1(\layer1[3][4] ), .ip2(n550), .ip3(reset), 
        .ip4(n549), .op(N1015) );
  nand2_1 U1087 ( .ip1(\layer1[2][4] ), .ip2(\layer1[3][4] ), .op(n553) );
  or2_1 U1088 ( .ip1(\layer1[2][4] ), .ip2(\layer1[3][4] ), .op(n551) );
  nand3_1 U1089 ( .ip1(\layer1[2][3] ), .ip2(\layer1[3][3] ), .ip3(n551), .op(
        n552) );
  nand2_1 U1090 ( .ip1(n553), .ip2(n552), .op(n555) );
  and2_1 U1091 ( .ip1(n554), .ip2(n778), .op(N1016) );
  fulladder U1092 ( .a(\layer1[2][5] ), .b(\layer1[3][5] ), .ci(n555), .co(
        n557), .s(n554) );
  and2_1 U1093 ( .ip1(n556), .ip2(n778), .op(N1017) );
  fulladder U1094 ( .a(\layer1[2][6] ), .b(\layer1[3][6] ), .ci(n557), .co(
        n559), .s(n556) );
  and2_1 U1095 ( .ip1(n558), .ip2(n672), .op(N1018) );
  fulladder U1096 ( .a(\layer1[2][7] ), .b(\layer1[3][7] ), .ci(n559), .co(
        n561), .s(n558) );
  and2_1 U1097 ( .ip1(n560), .ip2(n801), .op(N1019) );
  fulladder U1098 ( .a(\layer1[2][8] ), .b(\layer1[3][8] ), .ci(n561), .co(
        n563), .s(n560) );
  and2_1 U1099 ( .ip1(n562), .ip2(n672), .op(N1020) );
  fulladder U1100 ( .a(\layer1[2][9] ), .b(\layer1[3][9] ), .ci(n563), .co(
        n565), .s(n562) );
  and2_1 U1101 ( .ip1(n564), .ip2(n778), .op(N1021) );
  fulladder U1102 ( .a(\layer1[2][10] ), .b(\layer1[3][10] ), .ci(n565), .co(
        n567), .s(n564) );
  and2_1 U1103 ( .ip1(n566), .ip2(n672), .op(N1022) );
  fulladder U1104 ( .a(\layer1[2][11] ), .b(\layer1[3][11] ), .ci(n567), .co(
        n569), .s(n566) );
  and2_1 U1105 ( .ip1(n568), .ip2(n801), .op(N1023) );
  fulladder U1106 ( .a(\layer1[2][12] ), .b(\layer1[3][12] ), .ci(n569), .co(
        n571), .s(n568) );
  and2_1 U1107 ( .ip1(n570), .ip2(n801), .op(N1024) );
  fulladder U1108 ( .a(\layer1[2][13] ), .b(\layer1[3][13] ), .ci(n571), .co(
        n573), .s(n570) );
  and2_1 U1109 ( .ip1(n572), .ip2(n778), .op(N1025) );
  fulladder U1110 ( .a(\layer1[2][14] ), .b(\layer1[3][14] ), .ci(n573), .co(
        n575), .s(n572) );
  and2_1 U1111 ( .ip1(n574), .ip2(n672), .op(N1026) );
  fulladder U1112 ( .a(\layer1[2][15] ), .b(\layer1[3][15] ), .ci(n575), .co(
        n577), .s(n574) );
  and2_1 U1113 ( .ip1(n576), .ip2(n801), .op(N1027) );
  fulladder U1114 ( .a(\layer1[2][16] ), .b(\layer1[3][16] ), .ci(n577), .co(
        n579), .s(n576) );
  inv_1 U1115 ( .ip(reset), .op(n672) );
  and2_1 U1116 ( .ip1(n578), .ip2(n672), .op(N1028) );
  fulladder U1117 ( .a(\layer1[2][17] ), .b(\layer1[3][17] ), .ci(n579), .co(
        n581), .s(n578) );
  nor2_1 U1118 ( .ip1(n581), .ip2(\layer1[3][18] ), .op(n580) );
  not_ab_or_c_or_d U1119 ( .ip1(n581), .ip2(\layer1[3][18] ), .ip3(reset), 
        .ip4(n580), .op(N1029) );
  and3_1 U1120 ( .ip1(n581), .ip2(\layer1[3][18] ), .ip3(n801), .op(N1030) );
  and2_1 U1121 ( .ip1(N327), .ip2(n672), .op(N1047) );
  nor2_1 U1122 ( .ip1(\layer1[5][5] ), .ip2(\layer1[4][5] ), .op(n582) );
  nand2_1 U1123 ( .ip1(\layer1[5][5] ), .ip2(\layer1[4][5] ), .op(n583) );
  inv_1 U1124 ( .ip(n583), .op(n584) );
  nor3_1 U1125 ( .ip1(n582), .ip2(n483), .ip3(n584), .op(N1048) );
  mux2_1 U1126 ( .ip1(n584), .ip2(n583), .s(\layer1[4][6] ), .op(n586) );
  nor2_1 U1127 ( .ip1(\layer1[5][6] ), .ip2(n586), .op(n585) );
  not_ab_or_c_or_d U1128 ( .ip1(\layer1[5][6] ), .ip2(n586), .ip3(reset), 
        .ip4(n585), .op(N1049) );
  nand2_1 U1129 ( .ip1(\layer1[4][6] ), .ip2(\layer1[5][6] ), .op(n589) );
  or2_1 U1130 ( .ip1(\layer1[4][6] ), .ip2(\layer1[5][6] ), .op(n587) );
  nand3_1 U1131 ( .ip1(\layer1[4][5] ), .ip2(\layer1[5][5] ), .ip3(n587), .op(
        n588) );
  nand2_1 U1132 ( .ip1(n589), .ip2(n588), .op(n591) );
  and2_1 U1133 ( .ip1(n590), .ip2(n672), .op(N1050) );
  fulladder U1134 ( .a(\layer1[4][7] ), .b(\layer1[5][7] ), .ci(n591), .co(
        n593), .s(n590) );
  and2_1 U1135 ( .ip1(n592), .ip2(n672), .op(N1051) );
  fulladder U1136 ( .a(\layer1[4][8] ), .b(\layer1[5][8] ), .ci(n593), .co(
        n595), .s(n592) );
  and2_1 U1137 ( .ip1(n594), .ip2(n672), .op(N1052) );
  fulladder U1138 ( .a(\layer1[4][9] ), .b(\layer1[5][9] ), .ci(n595), .co(
        n597), .s(n594) );
  and2_1 U1139 ( .ip1(n596), .ip2(n672), .op(N1053) );
  fulladder U1140 ( .a(\layer1[4][10] ), .b(\layer1[5][10] ), .ci(n597), .co(
        n599), .s(n596) );
  and2_1 U1141 ( .ip1(n598), .ip2(n672), .op(N1054) );
  fulladder U1142 ( .a(\layer1[4][11] ), .b(\layer1[5][11] ), .ci(n599), .co(
        n601), .s(n598) );
  and2_1 U1143 ( .ip1(n600), .ip2(n672), .op(N1055) );
  fulladder U1144 ( .a(\layer1[4][12] ), .b(\layer1[5][12] ), .ci(n601), .co(
        n603), .s(n600) );
  and2_1 U1145 ( .ip1(n602), .ip2(n672), .op(N1056) );
  fulladder U1146 ( .a(\layer1[4][13] ), .b(\layer1[5][13] ), .ci(n603), .co(
        n605), .s(n602) );
  and2_1 U1147 ( .ip1(n604), .ip2(n672), .op(N1057) );
  fulladder U1148 ( .a(\layer1[4][14] ), .b(\layer1[5][14] ), .ci(n605), .co(
        n607), .s(n604) );
  and2_1 U1149 ( .ip1(n606), .ip2(n672), .op(N1058) );
  fulladder U1150 ( .a(\layer1[4][15] ), .b(\layer1[5][15] ), .ci(n607), .co(
        n609), .s(n606) );
  and2_1 U1151 ( .ip1(n608), .ip2(n672), .op(N1059) );
  fulladder U1152 ( .a(\layer1[4][16] ), .b(\layer1[5][16] ), .ci(n609), .co(
        n611), .s(n608) );
  and2_1 U1153 ( .ip1(n610), .ip2(n835), .op(N1060) );
  fulladder U1154 ( .a(\layer1[4][17] ), .b(\layer1[5][17] ), .ci(n611), .co(
        n613), .s(n610) );
  and2_1 U1155 ( .ip1(n612), .ip2(n835), .op(N1061) );
  fulladder U1156 ( .a(\layer1[4][18] ), .b(\layer1[5][18] ), .ci(n613), .co(
        n615), .s(n612) );
  and2_1 U1157 ( .ip1(n614), .ip2(n835), .op(N1062) );
  fulladder U1158 ( .a(\layer1[4][19] ), .b(\layer1[5][19] ), .ci(n615), .co(
        n617), .s(n614) );
  nor2_1 U1159 ( .ip1(n617), .ip2(\layer1[5][20] ), .op(n616) );
  not_ab_or_c_or_d U1160 ( .ip1(n617), .ip2(\layer1[5][20] ), .ip3(reset), 
        .ip4(n616), .op(N1063) );
  and3_1 U1161 ( .ip1(n617), .ip2(\layer1[5][20] ), .ip3(n835), .op(N1064) );
  and2_1 U1162 ( .ip1(N361), .ip2(n835), .op(N1081) );
  nor2_1 U1163 ( .ip1(\layer1[7][7] ), .ip2(\layer1[6][7] ), .op(n618) );
  nand2_1 U1164 ( .ip1(\layer1[7][7] ), .ip2(\layer1[6][7] ), .op(n619) );
  inv_1 U1165 ( .ip(n619), .op(n620) );
  nor3_1 U1166 ( .ip1(n618), .ip2(n483), .ip3(n620), .op(N1082) );
  mux2_1 U1167 ( .ip1(n620), .ip2(n619), .s(\layer1[6][8] ), .op(n622) );
  nor2_1 U1168 ( .ip1(\layer1[7][8] ), .ip2(n622), .op(n621) );
  not_ab_or_c_or_d U1169 ( .ip1(\layer1[7][8] ), .ip2(n622), .ip3(reset), 
        .ip4(n621), .op(N1083) );
  nand2_1 U1170 ( .ip1(\layer1[6][8] ), .ip2(\layer1[7][8] ), .op(n625) );
  or2_1 U1171 ( .ip1(\layer1[6][8] ), .ip2(\layer1[7][8] ), .op(n623) );
  nand3_1 U1172 ( .ip1(\layer1[6][7] ), .ip2(\layer1[7][7] ), .ip3(n623), .op(
        n624) );
  nand2_1 U1173 ( .ip1(n625), .ip2(n624), .op(n627) );
  and2_1 U1174 ( .ip1(n626), .ip2(n835), .op(N1084) );
  fulladder U1175 ( .a(\layer1[6][9] ), .b(\layer1[7][9] ), .ci(n627), .co(
        n629), .s(n626) );
  and2_1 U1176 ( .ip1(n628), .ip2(n835), .op(N1085) );
  fulladder U1177 ( .a(\layer1[6][10] ), .b(\layer1[7][10] ), .ci(n629), .co(
        n631), .s(n628) );
  and2_1 U1178 ( .ip1(n630), .ip2(n835), .op(N1086) );
  fulladder U1179 ( .a(\layer1[6][11] ), .b(\layer1[7][11] ), .ci(n631), .co(
        n633), .s(n630) );
  and2_1 U1180 ( .ip1(n632), .ip2(n835), .op(N1087) );
  fulladder U1181 ( .a(\layer1[6][12] ), .b(\layer1[7][12] ), .ci(n633), .co(
        n635), .s(n632) );
  and2_1 U1182 ( .ip1(n634), .ip2(n835), .op(N1088) );
  fulladder U1183 ( .a(\layer1[6][13] ), .b(\layer1[7][13] ), .ci(n635), .co(
        n637), .s(n634) );
  and2_1 U1184 ( .ip1(n636), .ip2(n835), .op(N1089) );
  fulladder U1185 ( .a(\layer1[6][14] ), .b(\layer1[7][14] ), .ci(n637), .co(
        n639), .s(n636) );
  and2_1 U1186 ( .ip1(n638), .ip2(n835), .op(N1090) );
  fulladder U1187 ( .a(\layer1[6][15] ), .b(\layer1[7][15] ), .ci(n639), .co(
        n641), .s(n638) );
  and2_1 U1188 ( .ip1(n640), .ip2(n835), .op(N1091) );
  fulladder U1189 ( .a(\layer1[6][16] ), .b(\layer1[7][16] ), .ci(n641), .co(
        n643), .s(n640) );
  and2_1 U1190 ( .ip1(n642), .ip2(n672), .op(N1092) );
  fulladder U1191 ( .a(\layer1[6][17] ), .b(\layer1[7][17] ), .ci(n643), .co(
        n645), .s(n642) );
  and2_1 U1192 ( .ip1(n644), .ip2(n672), .op(N1093) );
  fulladder U1193 ( .a(\layer1[6][18] ), .b(\layer1[7][18] ), .ci(n645), .co(
        n647), .s(n644) );
  and2_1 U1194 ( .ip1(n646), .ip2(n672), .op(N1094) );
  fulladder U1195 ( .a(\layer1[6][19] ), .b(\layer1[7][19] ), .ci(n647), .co(
        n649), .s(n646) );
  and2_1 U1196 ( .ip1(n648), .ip2(n672), .op(N1095) );
  fulladder U1197 ( .a(\layer1[6][20] ), .b(\layer1[7][20] ), .ci(n649), .co(
        n651), .s(n648) );
  and2_1 U1198 ( .ip1(n650), .ip2(n672), .op(N1096) );
  fulladder U1199 ( .a(\layer1[6][21] ), .b(\layer1[7][21] ), .ci(n651), .co(
        n653), .s(n650) );
  nor2_1 U1200 ( .ip1(n653), .ip2(\layer1[7][22] ), .op(n652) );
  not_ab_or_c_or_d U1201 ( .ip1(n653), .ip2(\layer1[7][22] ), .ip3(reset), 
        .ip4(n652), .op(N1097) );
  and3_1 U1202 ( .ip1(n653), .ip2(\layer1[7][22] ), .ip3(n801), .op(N1098) );
  and2_1 U1203 ( .ip1(N395), .ip2(n672), .op(N1115) );
  nor2_1 U1204 ( .ip1(\layer1[9][9] ), .ip2(\layer1[8][9] ), .op(n654) );
  nand2_1 U1205 ( .ip1(\layer1[9][9] ), .ip2(\layer1[8][9] ), .op(n655) );
  inv_1 U1206 ( .ip(n655), .op(n656) );
  nor3_1 U1207 ( .ip1(n654), .ip2(n483), .ip3(n656), .op(N1116) );
  mux2_1 U1208 ( .ip1(n656), .ip2(n655), .s(\layer1[8][10] ), .op(n658) );
  nor2_1 U1209 ( .ip1(\layer1[9][10] ), .ip2(n658), .op(n657) );
  not_ab_or_c_or_d U1210 ( .ip1(\layer1[9][10] ), .ip2(n658), .ip3(reset), 
        .ip4(n657), .op(N1117) );
  nand2_1 U1211 ( .ip1(\layer1[8][10] ), .ip2(\layer1[9][10] ), .op(n661) );
  or2_1 U1212 ( .ip1(\layer1[8][10] ), .ip2(\layer1[9][10] ), .op(n659) );
  nand3_1 U1213 ( .ip1(\layer1[8][9] ), .ip2(\layer1[9][9] ), .ip3(n659), .op(
        n660) );
  nand2_1 U1214 ( .ip1(n661), .ip2(n660), .op(n663) );
  and2_1 U1215 ( .ip1(n662), .ip2(n672), .op(N1118) );
  fulladder U1216 ( .a(\layer1[8][11] ), .b(\layer1[9][11] ), .ci(n663), .co(
        n665), .s(n662) );
  and2_1 U1217 ( .ip1(n664), .ip2(n672), .op(N1119) );
  fulladder U1218 ( .a(\layer1[8][12] ), .b(\layer1[9][12] ), .ci(n665), .co(
        n667), .s(n664) );
  and2_1 U1219 ( .ip1(n666), .ip2(n672), .op(N1120) );
  fulladder U1220 ( .a(\layer1[8][13] ), .b(\layer1[9][13] ), .ci(n667), .co(
        n669), .s(n666) );
  and2_1 U1221 ( .ip1(n668), .ip2(n672), .op(N1121) );
  fulladder U1222 ( .a(\layer1[8][14] ), .b(\layer1[9][14] ), .ci(n669), .co(
        n671), .s(n668) );
  and2_1 U1223 ( .ip1(n670), .ip2(n672), .op(N1122) );
  fulladder U1224 ( .a(\layer1[8][15] ), .b(\layer1[9][15] ), .ci(n671), .co(
        n674), .s(n670) );
  and2_1 U1225 ( .ip1(n673), .ip2(n672), .op(N1123) );
  fulladder U1226 ( .a(\layer1[8][16] ), .b(\layer1[9][16] ), .ci(n674), .co(
        n676), .s(n673) );
  and2_1 U1227 ( .ip1(n675), .ip2(n540), .op(N1124) );
  fulladder U1228 ( .a(\layer1[8][17] ), .b(\layer1[9][17] ), .ci(n676), .co(
        n678), .s(n675) );
  and2_1 U1229 ( .ip1(n677), .ip2(n672), .op(N1125) );
  fulladder U1230 ( .a(\layer1[8][18] ), .b(\layer1[9][18] ), .ci(n678), .co(
        n680), .s(n677) );
  and2_1 U1231 ( .ip1(n679), .ip2(n801), .op(N1126) );
  fulladder U1232 ( .a(\layer1[8][19] ), .b(\layer1[9][19] ), .ci(n680), .co(
        n682), .s(n679) );
  and2_1 U1233 ( .ip1(n681), .ip2(n778), .op(N1127) );
  fulladder U1234 ( .a(\layer1[8][20] ), .b(\layer1[9][20] ), .ci(n682), .co(
        n684), .s(n681) );
  and2_1 U1235 ( .ip1(n683), .ip2(n835), .op(N1128) );
  fulladder U1236 ( .a(\layer1[8][21] ), .b(\layer1[9][21] ), .ci(n684), .co(
        n686), .s(n683) );
  and2_1 U1237 ( .ip1(n685), .ip2(n540), .op(N1129) );
  fulladder U1238 ( .a(\layer1[8][22] ), .b(\layer1[9][22] ), .ci(n686), .co(
        n688), .s(n685) );
  xor2_1 U1239 ( .ip1(\layer1[9][23] ), .ip2(\layer1[8][23] ), .op(n687) );
  xor2_1 U1240 ( .ip1(n688), .ip2(n687), .op(n689) );
  and2_1 U1241 ( .ip1(n689), .ip2(n672), .op(N1130) );
  and2_1 U1242 ( .ip1(N429), .ip2(n801), .op(N1149) );
  nor2_1 U1243 ( .ip1(\layer1[11][11] ), .ip2(\layer1[10][11] ), .op(n690) );
  nand2_1 U1244 ( .ip1(\layer1[11][11] ), .ip2(\layer1[10][11] ), .op(n691) );
  inv_1 U1245 ( .ip(n691), .op(n692) );
  nor3_1 U1246 ( .ip1(n690), .ip2(n483), .ip3(n692), .op(N1150) );
  mux2_1 U1247 ( .ip1(n692), .ip2(n691), .s(\layer1[10][12] ), .op(n694) );
  nor2_1 U1248 ( .ip1(\layer1[11][12] ), .ip2(n694), .op(n693) );
  not_ab_or_c_or_d U1249 ( .ip1(\layer1[11][12] ), .ip2(n694), .ip3(reset), 
        .ip4(n693), .op(N1151) );
  nand2_1 U1250 ( .ip1(\layer1[10][12] ), .ip2(\layer1[11][12] ), .op(n697) );
  or2_1 U1251 ( .ip1(\layer1[10][12] ), .ip2(\layer1[11][12] ), .op(n695) );
  nand3_1 U1252 ( .ip1(\layer1[10][11] ), .ip2(\layer1[11][11] ), .ip3(n695), 
        .op(n696) );
  nand2_1 U1253 ( .ip1(n697), .ip2(n696), .op(n699) );
  and2_1 U1254 ( .ip1(n698), .ip2(n778), .op(N1152) );
  fulladder U1255 ( .a(\layer1[10][13] ), .b(\layer1[11][13] ), .ci(n699), 
        .co(n701), .s(n698) );
  and2_1 U1256 ( .ip1(n700), .ip2(n835), .op(N1153) );
  fulladder U1257 ( .a(\layer1[10][14] ), .b(\layer1[11][14] ), .ci(n701), 
        .co(n703), .s(n700) );
  and2_1 U1258 ( .ip1(n702), .ip2(n540), .op(N1154) );
  fulladder U1259 ( .a(\layer1[10][15] ), .b(\layer1[11][15] ), .ci(n703), 
        .co(n705), .s(n702) );
  and2_1 U1260 ( .ip1(n704), .ip2(n672), .op(N1155) );
  fulladder U1261 ( .a(\layer1[10][16] ), .b(\layer1[11][16] ), .ci(n705), 
        .co(n707), .s(n704) );
  and2_1 U1262 ( .ip1(n706), .ip2(n801), .op(N1156) );
  fulladder U1263 ( .a(\layer1[10][17] ), .b(\layer1[11][17] ), .ci(n707), 
        .co(n709), .s(n706) );
  and2_1 U1264 ( .ip1(n708), .ip2(n778), .op(N1157) );
  fulladder U1265 ( .a(\layer1[10][18] ), .b(\layer1[11][18] ), .ci(n709), 
        .co(n711), .s(n708) );
  and2_1 U1266 ( .ip1(n710), .ip2(n835), .op(N1158) );
  fulladder U1267 ( .a(\layer1[10][19] ), .b(\layer1[11][19] ), .ci(n711), 
        .co(n713), .s(n710) );
  and2_1 U1268 ( .ip1(n712), .ip2(n540), .op(N1159) );
  fulladder U1269 ( .a(\layer1[10][20] ), .b(\layer1[11][20] ), .ci(n713), 
        .co(n715), .s(n712) );
  and2_1 U1270 ( .ip1(n714), .ip2(n672), .op(N1160) );
  fulladder U1271 ( .a(\layer1[10][21] ), .b(\layer1[11][21] ), .ci(n715), 
        .co(n717), .s(n714) );
  and2_1 U1272 ( .ip1(n716), .ip2(n801), .op(N1161) );
  fulladder U1273 ( .a(\layer1[10][22] ), .b(\layer1[11][22] ), .ci(n717), 
        .co(n719), .s(n716) );
  xor2_1 U1274 ( .ip1(\layer1[11][23] ), .ip2(\layer1[10][23] ), .op(n718) );
  xor2_1 U1275 ( .ip1(n719), .ip2(n718), .op(n720) );
  and2_1 U1276 ( .ip1(n720), .ip2(n778), .op(N1162) );
  and2_1 U1277 ( .ip1(N463), .ip2(n835), .op(N1183) );
  nor2_1 U1278 ( .ip1(\layer1[13][13] ), .ip2(\layer1[12][13] ), .op(n721) );
  nand2_1 U1279 ( .ip1(\layer1[13][13] ), .ip2(\layer1[12][13] ), .op(n722) );
  inv_1 U1280 ( .ip(n722), .op(n723) );
  nor3_1 U1281 ( .ip1(n721), .ip2(n483), .ip3(n723), .op(N1184) );
  mux2_1 U1282 ( .ip1(n723), .ip2(n722), .s(\layer1[12][14] ), .op(n725) );
  nor2_1 U1283 ( .ip1(\layer1[13][14] ), .ip2(n725), .op(n724) );
  not_ab_or_c_or_d U1284 ( .ip1(\layer1[13][14] ), .ip2(n725), .ip3(reset), 
        .ip4(n724), .op(N1185) );
  nand2_1 U1285 ( .ip1(\layer1[12][14] ), .ip2(\layer1[13][14] ), .op(n728) );
  or2_1 U1286 ( .ip1(\layer1[12][14] ), .ip2(\layer1[13][14] ), .op(n726) );
  nand3_1 U1287 ( .ip1(\layer1[12][13] ), .ip2(\layer1[13][13] ), .ip3(n726), 
        .op(n727) );
  nand2_1 U1288 ( .ip1(n728), .ip2(n727), .op(n730) );
  and2_1 U1289 ( .ip1(n729), .ip2(n540), .op(N1186) );
  fulladder U1290 ( .a(\layer1[12][15] ), .b(\layer1[13][15] ), .ci(n730), 
        .co(n732), .s(n729) );
  and2_1 U1291 ( .ip1(n731), .ip2(n672), .op(N1187) );
  fulladder U1292 ( .a(\layer1[12][16] ), .b(\layer1[13][16] ), .ci(n732), 
        .co(n734), .s(n731) );
  and2_1 U1293 ( .ip1(n733), .ip2(n801), .op(N1188) );
  fulladder U1294 ( .a(\layer1[12][17] ), .b(\layer1[13][17] ), .ci(n734), 
        .co(n736), .s(n733) );
  and2_1 U1295 ( .ip1(n735), .ip2(n778), .op(N1189) );
  fulladder U1296 ( .a(\layer1[12][18] ), .b(\layer1[13][18] ), .ci(n736), 
        .co(n738), .s(n735) );
  and2_1 U1297 ( .ip1(n737), .ip2(n778), .op(N1190) );
  fulladder U1298 ( .a(\layer1[12][19] ), .b(\layer1[13][19] ), .ci(n738), 
        .co(n740), .s(n737) );
  and2_1 U1299 ( .ip1(n739), .ip2(n778), .op(N1191) );
  fulladder U1300 ( .a(\layer1[12][20] ), .b(\layer1[13][20] ), .ci(n740), 
        .co(n742), .s(n739) );
  and2_1 U1301 ( .ip1(n741), .ip2(n672), .op(N1192) );
  fulladder U1302 ( .a(\layer1[12][21] ), .b(\layer1[13][21] ), .ci(n742), 
        .co(n744), .s(n741) );
  and2_1 U1303 ( .ip1(n743), .ip2(n801), .op(N1193) );
  fulladder U1304 ( .a(\layer1[12][22] ), .b(\layer1[13][22] ), .ci(n744), 
        .co(n747), .s(n743) );
  xor2_1 U1305 ( .ip1(\layer1[13][23] ), .ip2(\layer1[12][23] ), .op(n746) );
  nor2_1 U1306 ( .ip1(n747), .ip2(n746), .op(n745) );
  not_ab_or_c_or_d U1307 ( .ip1(n747), .ip2(n746), .ip3(reset), .ip4(n745), 
        .op(N1194) );
  and2_1 U1308 ( .ip1(N497), .ip2(n672), .op(N1217) );
  nor2_1 U1309 ( .ip1(\layer1[15][15] ), .ip2(\layer1[14][15] ), .op(n748) );
  nand2_1 U1310 ( .ip1(\layer1[15][15] ), .ip2(\layer1[14][15] ), .op(n749) );
  inv_1 U1311 ( .ip(n749), .op(n750) );
  nor3_1 U1312 ( .ip1(n748), .ip2(n483), .ip3(n750), .op(N1218) );
  mux2_1 U1313 ( .ip1(n750), .ip2(n749), .s(\layer1[14][16] ), .op(n752) );
  nor2_1 U1314 ( .ip1(\layer1[15][16] ), .ip2(n752), .op(n751) );
  not_ab_or_c_or_d U1315 ( .ip1(\layer1[15][16] ), .ip2(n752), .ip3(reset), 
        .ip4(n751), .op(N1219) );
  nand2_1 U1316 ( .ip1(\layer1[14][16] ), .ip2(\layer1[15][16] ), .op(n755) );
  or2_1 U1317 ( .ip1(\layer1[14][16] ), .ip2(\layer1[15][16] ), .op(n753) );
  nand3_1 U1318 ( .ip1(\layer1[14][15] ), .ip2(\layer1[15][15] ), .ip3(n753), 
        .op(n754) );
  nand2_1 U1319 ( .ip1(n755), .ip2(n754), .op(n757) );
  and2_1 U1320 ( .ip1(n756), .ip2(n778), .op(N1220) );
  fulladder U1321 ( .a(\layer1[14][17] ), .b(\layer1[15][17] ), .ci(n757), 
        .co(n759), .s(n756) );
  and2_1 U1322 ( .ip1(n758), .ip2(n672), .op(N1221) );
  fulladder U1323 ( .a(\layer1[14][18] ), .b(\layer1[15][18] ), .ci(n759), 
        .co(n761), .s(n758) );
  and2_1 U1324 ( .ip1(n760), .ip2(n801), .op(N1222) );
  fulladder U1325 ( .a(\layer1[14][19] ), .b(\layer1[15][19] ), .ci(n761), 
        .co(n763), .s(n760) );
  and2_1 U1326 ( .ip1(n762), .ip2(n801), .op(N1223) );
  fulladder U1327 ( .a(\layer1[14][20] ), .b(\layer1[15][20] ), .ci(n763), 
        .co(n765), .s(n762) );
  and2_1 U1328 ( .ip1(n764), .ip2(n778), .op(N1224) );
  fulladder U1329 ( .a(\layer1[14][21] ), .b(\layer1[15][21] ), .ci(n765), 
        .co(n767), .s(n764) );
  and2_1 U1330 ( .ip1(n766), .ip2(n672), .op(N1225) );
  fulladder U1331 ( .a(\layer1[14][22] ), .b(\layer1[15][22] ), .ci(n767), 
        .co(n770), .s(n766) );
  xor2_1 U1332 ( .ip1(\layer1[15][23] ), .ip2(\layer1[14][23] ), .op(n769) );
  nor2_1 U1333 ( .ip1(n770), .ip2(n769), .op(n768) );
  not_ab_or_c_or_d U1334 ( .ip1(n770), .ip2(n769), .ip3(reset), .ip4(n768), 
        .op(N1226) );
  inv_1 U1335 ( .ip(in[1]), .op(n787) );
  nand2_1 U1336 ( .ip1(w[0]), .ip2(n801), .op(n771) );
  nor2_1 U1337 ( .ip1(n787), .ip2(n771), .op(N724) );
  inv_1 U1338 ( .ip(in[2]), .op(n788) );
  nor2_1 U1339 ( .ip1(n788), .ip2(n771), .op(N725) );
  inv_1 U1340 ( .ip(in[3]), .op(n789) );
  nor2_1 U1341 ( .ip1(n789), .ip2(n771), .op(N726) );
  inv_1 U1342 ( .ip(in[4]), .op(n790) );
  nor2_1 U1343 ( .ip1(n790), .ip2(n771), .op(N727) );
  inv_1 U1344 ( .ip(in[5]), .op(n791) );
  nor2_1 U1345 ( .ip1(n791), .ip2(n771), .op(N728) );
  inv_1 U1346 ( .ip(in[6]), .op(n792) );
  nor2_1 U1347 ( .ip1(n792), .ip2(n771), .op(N729) );
  inv_1 U1348 ( .ip(in[7]), .op(n793) );
  nor2_1 U1349 ( .ip1(n793), .ip2(n771), .op(N730) );
  inv_1 U1350 ( .ip(in[8]), .op(n794) );
  nor2_1 U1351 ( .ip1(n794), .ip2(n771), .op(N731) );
  inv_1 U1352 ( .ip(in[9]), .op(n795) );
  nor2_1 U1353 ( .ip1(n771), .ip2(n795), .op(N732) );
  inv_1 U1354 ( .ip(in[10]), .op(n800) );
  nor2_1 U1355 ( .ip1(n771), .ip2(n800), .op(N733) );
  inv_1 U1356 ( .ip(in[11]), .op(n797) );
  nor2_1 U1357 ( .ip1(n771), .ip2(n797), .op(N734) );
  inv_1 U1358 ( .ip(in[12]), .op(n781) );
  nor2_1 U1359 ( .ip1(n771), .ip2(n781), .op(N735) );
  inv_1 U1360 ( .ip(in[13]), .op(n785) );
  nor2_1 U1361 ( .ip1(n771), .ip2(n785), .op(N736) );
  inv_1 U1362 ( .ip(in[14]), .op(n783) );
  nor2_1 U1363 ( .ip1(n771), .ip2(n783), .op(N737) );
  inv_1 U1364 ( .ip(in[0]), .op(n798) );
  nand2_1 U1365 ( .ip1(w[1]), .ip2(n778), .op(n772) );
  nor2_1 U1366 ( .ip1(n798), .ip2(n772), .op(N739) );
  nor2_1 U1367 ( .ip1(n787), .ip2(n772), .op(N740) );
  nor2_1 U1368 ( .ip1(n788), .ip2(n772), .op(N741) );
  nor2_1 U1369 ( .ip1(n789), .ip2(n772), .op(N742) );
  nor2_1 U1370 ( .ip1(n790), .ip2(n772), .op(N743) );
  nor2_1 U1371 ( .ip1(n791), .ip2(n772), .op(N744) );
  nor2_1 U1372 ( .ip1(n792), .ip2(n772), .op(N745) );
  nor2_1 U1373 ( .ip1(n793), .ip2(n772), .op(N746) );
  nor2_1 U1374 ( .ip1(n794), .ip2(n772), .op(N747) );
  nor2_1 U1375 ( .ip1(n795), .ip2(n772), .op(N748) );
  nor2_1 U1376 ( .ip1(n800), .ip2(n772), .op(N749) );
  nor2_1 U1377 ( .ip1(n797), .ip2(n772), .op(N750) );
  nor2_1 U1378 ( .ip1(n781), .ip2(n772), .op(N751) );
  nor2_1 U1379 ( .ip1(n785), .ip2(n772), .op(N752) );
  nor2_1 U1380 ( .ip1(n783), .ip2(n772), .op(N753) );
  nand2_1 U1381 ( .ip1(w[2]), .ip2(n801), .op(n773) );
  nor2_1 U1382 ( .ip1(n798), .ip2(n773), .op(N755) );
  nor2_1 U1383 ( .ip1(n787), .ip2(n773), .op(N756) );
  nor2_1 U1384 ( .ip1(n788), .ip2(n773), .op(N757) );
  nor2_1 U1385 ( .ip1(n789), .ip2(n773), .op(N758) );
  nor2_1 U1386 ( .ip1(n790), .ip2(n773), .op(N759) );
  nor2_1 U1387 ( .ip1(n791), .ip2(n773), .op(N760) );
  nor2_1 U1388 ( .ip1(n792), .ip2(n773), .op(N761) );
  nor2_1 U1389 ( .ip1(n793), .ip2(n773), .op(N762) );
  nor2_1 U1390 ( .ip1(n794), .ip2(n773), .op(N763) );
  nor2_1 U1391 ( .ip1(n795), .ip2(n773), .op(N764) );
  nor2_1 U1392 ( .ip1(n800), .ip2(n773), .op(N765) );
  nor2_1 U1393 ( .ip1(n797), .ip2(n773), .op(N766) );
  nor2_1 U1394 ( .ip1(n781), .ip2(n773), .op(N767) );
  nor2_1 U1395 ( .ip1(n785), .ip2(n773), .op(N768) );
  nor2_1 U1396 ( .ip1(n783), .ip2(n773), .op(N769) );
  nand2_1 U1397 ( .ip1(w[3]), .ip2(n801), .op(n774) );
  nor2_1 U1398 ( .ip1(n798), .ip2(n774), .op(N771) );
  nor2_1 U1399 ( .ip1(n787), .ip2(n774), .op(N772) );
  nor2_1 U1400 ( .ip1(n788), .ip2(n774), .op(N773) );
  nor2_1 U1401 ( .ip1(n789), .ip2(n774), .op(N774) );
  nor2_1 U1402 ( .ip1(n790), .ip2(n774), .op(N775) );
  nor2_1 U1403 ( .ip1(n791), .ip2(n774), .op(N776) );
  nor2_1 U1404 ( .ip1(n792), .ip2(n774), .op(N777) );
  nor2_1 U1405 ( .ip1(n793), .ip2(n774), .op(N778) );
  nor2_1 U1406 ( .ip1(n794), .ip2(n774), .op(N779) );
  nor2_1 U1407 ( .ip1(n795), .ip2(n774), .op(N780) );
  nor2_1 U1408 ( .ip1(n800), .ip2(n774), .op(N781) );
  nor2_1 U1409 ( .ip1(n797), .ip2(n774), .op(N782) );
  nor2_1 U1410 ( .ip1(n781), .ip2(n774), .op(N783) );
  nor2_1 U1411 ( .ip1(n785), .ip2(n774), .op(N784) );
  nor2_1 U1412 ( .ip1(n783), .ip2(n774), .op(N785) );
  nand2_1 U1413 ( .ip1(w[4]), .ip2(n801), .op(n775) );
  nor2_1 U1414 ( .ip1(n798), .ip2(n775), .op(N787) );
  nor2_1 U1415 ( .ip1(n787), .ip2(n775), .op(N788) );
  nor2_1 U1416 ( .ip1(n788), .ip2(n775), .op(N789) );
  nor2_1 U1417 ( .ip1(n789), .ip2(n775), .op(N790) );
  nor2_1 U1418 ( .ip1(n790), .ip2(n775), .op(N791) );
  nor2_1 U1419 ( .ip1(n791), .ip2(n775), .op(N792) );
  nor2_1 U1420 ( .ip1(n792), .ip2(n775), .op(N793) );
  nor2_1 U1421 ( .ip1(n793), .ip2(n775), .op(N794) );
  nor2_1 U1422 ( .ip1(n794), .ip2(n775), .op(N795) );
  nor2_1 U1423 ( .ip1(n795), .ip2(n775), .op(N796) );
  nor2_1 U1424 ( .ip1(n800), .ip2(n775), .op(N797) );
  nor2_1 U1425 ( .ip1(n797), .ip2(n775), .op(N798) );
  nor2_1 U1426 ( .ip1(n781), .ip2(n775), .op(N799) );
  nor2_1 U1427 ( .ip1(n785), .ip2(n775), .op(N800) );
  nor2_1 U1428 ( .ip1(n783), .ip2(n775), .op(N801) );
  nand2_1 U1429 ( .ip1(w[5]), .ip2(n778), .op(n776) );
  nor2_1 U1430 ( .ip1(n798), .ip2(n776), .op(N803) );
  nor2_1 U1431 ( .ip1(n787), .ip2(n776), .op(N804) );
  nor2_1 U1432 ( .ip1(n788), .ip2(n776), .op(N805) );
  nor2_1 U1433 ( .ip1(n789), .ip2(n776), .op(N806) );
  nor2_1 U1434 ( .ip1(n790), .ip2(n776), .op(N807) );
  nor2_1 U1435 ( .ip1(n791), .ip2(n776), .op(N808) );
  nor2_1 U1436 ( .ip1(n792), .ip2(n776), .op(N809) );
  nor2_1 U1437 ( .ip1(n793), .ip2(n776), .op(N810) );
  nor2_1 U1438 ( .ip1(n794), .ip2(n776), .op(N811) );
  nor2_1 U1439 ( .ip1(n795), .ip2(n776), .op(N812) );
  nor2_1 U1440 ( .ip1(n800), .ip2(n776), .op(N813) );
  nor2_1 U1441 ( .ip1(n797), .ip2(n776), .op(N814) );
  nor2_1 U1442 ( .ip1(n781), .ip2(n776), .op(N815) );
  nor2_1 U1443 ( .ip1(n785), .ip2(n776), .op(N816) );
  nor2_1 U1444 ( .ip1(n783), .ip2(n776), .op(N817) );
  nand2_1 U1445 ( .ip1(w[6]), .ip2(n801), .op(n777) );
  nor2_1 U1446 ( .ip1(n798), .ip2(n777), .op(N819) );
  nor2_1 U1447 ( .ip1(n787), .ip2(n777), .op(N820) );
  nor2_1 U1448 ( .ip1(n788), .ip2(n777), .op(N821) );
  nor2_1 U1449 ( .ip1(n789), .ip2(n777), .op(N822) );
  nor2_1 U1450 ( .ip1(n790), .ip2(n777), .op(N823) );
  nor2_1 U1451 ( .ip1(n791), .ip2(n777), .op(N824) );
  nor2_1 U1452 ( .ip1(n792), .ip2(n777), .op(N825) );
  nor2_1 U1453 ( .ip1(n793), .ip2(n777), .op(N826) );
  nor2_1 U1454 ( .ip1(n794), .ip2(n777), .op(N827) );
  nor2_1 U1455 ( .ip1(n795), .ip2(n777), .op(N828) );
  nor2_1 U1456 ( .ip1(n800), .ip2(n777), .op(N829) );
  nor2_1 U1457 ( .ip1(n797), .ip2(n777), .op(N830) );
  nor2_1 U1458 ( .ip1(n781), .ip2(n777), .op(N831) );
  nor2_1 U1459 ( .ip1(n785), .ip2(n777), .op(N832) );
  nor2_1 U1460 ( .ip1(n783), .ip2(n777), .op(N833) );
  nand2_1 U1461 ( .ip1(w[7]), .ip2(n778), .op(n779) );
  nor2_1 U1462 ( .ip1(n798), .ip2(n779), .op(N835) );
  nor2_1 U1463 ( .ip1(n787), .ip2(n779), .op(N836) );
  nor2_1 U1464 ( .ip1(n788), .ip2(n779), .op(N837) );
  nor2_1 U1465 ( .ip1(n789), .ip2(n779), .op(N838) );
  nor2_1 U1466 ( .ip1(n790), .ip2(n779), .op(N839) );
  nor2_1 U1467 ( .ip1(n791), .ip2(n779), .op(N840) );
  nor2_1 U1468 ( .ip1(n792), .ip2(n779), .op(N841) );
  nor2_1 U1469 ( .ip1(n793), .ip2(n779), .op(N842) );
  nor2_1 U1470 ( .ip1(n794), .ip2(n779), .op(N843) );
  nor2_1 U1471 ( .ip1(n795), .ip2(n779), .op(N844) );
  nor2_1 U1472 ( .ip1(n800), .ip2(n779), .op(N845) );
  nor2_1 U1473 ( .ip1(n797), .ip2(n779), .op(N846) );
  nor2_1 U1474 ( .ip1(n781), .ip2(n779), .op(N847) );
  nor2_1 U1475 ( .ip1(n785), .ip2(n779), .op(N848) );
  nor2_1 U1476 ( .ip1(n783), .ip2(n779), .op(N849) );
  nand2_1 U1477 ( .ip1(w[8]), .ip2(n801), .op(n780) );
  nor2_1 U1478 ( .ip1(n798), .ip2(n780), .op(N851) );
  nor2_1 U1479 ( .ip1(n787), .ip2(n780), .op(N852) );
  nor2_1 U1480 ( .ip1(n788), .ip2(n780), .op(N853) );
  nor2_1 U1481 ( .ip1(n789), .ip2(n780), .op(N854) );
  nor2_1 U1482 ( .ip1(n790), .ip2(n780), .op(N855) );
  nor2_1 U1483 ( .ip1(n791), .ip2(n780), .op(N856) );
  nor2_1 U1484 ( .ip1(n792), .ip2(n780), .op(N857) );
  nor2_1 U1485 ( .ip1(n793), .ip2(n780), .op(N858) );
  nor2_1 U1486 ( .ip1(n794), .ip2(n780), .op(N859) );
  nor2_1 U1487 ( .ip1(n795), .ip2(n780), .op(N860) );
  nor2_1 U1488 ( .ip1(n800), .ip2(n780), .op(N861) );
  nor2_1 U1489 ( .ip1(n797), .ip2(n780), .op(N862) );
  nor2_1 U1490 ( .ip1(n781), .ip2(n780), .op(N863) );
  nor2_1 U1491 ( .ip1(n785), .ip2(n780), .op(N864) );
  nor2_1 U1492 ( .ip1(n783), .ip2(n780), .op(N865) );
  nand2_1 U1493 ( .ip1(w[9]), .ip2(n801), .op(n782) );
  nor2_1 U1494 ( .ip1(n798), .ip2(n782), .op(N867) );
  nor2_1 U1495 ( .ip1(n787), .ip2(n782), .op(N868) );
  nor2_1 U1496 ( .ip1(n788), .ip2(n782), .op(N869) );
  nor2_1 U1497 ( .ip1(n789), .ip2(n782), .op(N870) );
  nor2_1 U1498 ( .ip1(n790), .ip2(n782), .op(N871) );
  nor2_1 U1499 ( .ip1(n791), .ip2(n782), .op(N872) );
  nor2_1 U1500 ( .ip1(n792), .ip2(n782), .op(N873) );
  nor2_1 U1501 ( .ip1(n793), .ip2(n782), .op(N874) );
  nor2_1 U1502 ( .ip1(n794), .ip2(n782), .op(N875) );
  nor2_1 U1503 ( .ip1(n795), .ip2(n782), .op(N876) );
  nor2_1 U1504 ( .ip1(n800), .ip2(n782), .op(N877) );
  nor2_1 U1505 ( .ip1(n797), .ip2(n782), .op(N878) );
  nor2_1 U1506 ( .ip1(n781), .ip2(n782), .op(N879) );
  nor2_1 U1507 ( .ip1(n785), .ip2(n782), .op(N880) );
  nor2_1 U1508 ( .ip1(n783), .ip2(n782), .op(N881) );
  nand2_1 U1509 ( .ip1(w[10]), .ip2(n801), .op(n784) );
  nor2_1 U1510 ( .ip1(n798), .ip2(n784), .op(N883) );
  nor2_1 U1511 ( .ip1(n787), .ip2(n784), .op(N884) );
  nor2_1 U1512 ( .ip1(n788), .ip2(n784), .op(N885) );
  nor2_1 U1513 ( .ip1(n789), .ip2(n784), .op(N886) );
  nor2_1 U1514 ( .ip1(n790), .ip2(n784), .op(N887) );
  nor2_1 U1515 ( .ip1(n791), .ip2(n784), .op(N888) );
  nor2_1 U1516 ( .ip1(n792), .ip2(n784), .op(N889) );
  nor2_1 U1517 ( .ip1(n793), .ip2(n784), .op(N890) );
  nor2_1 U1518 ( .ip1(n794), .ip2(n784), .op(N891) );
  nor2_1 U1519 ( .ip1(n795), .ip2(n784), .op(N892) );
  nor2_1 U1520 ( .ip1(n800), .ip2(n784), .op(N893) );
  nor2_1 U1521 ( .ip1(n797), .ip2(n784), .op(N894) );
  nor2_1 U1522 ( .ip1(n781), .ip2(n784), .op(N895) );
  nor2_1 U1523 ( .ip1(n785), .ip2(n784), .op(N896) );
  nand2_1 U1524 ( .ip1(w[11]), .ip2(n801), .op(n786) );
  nor2_1 U1525 ( .ip1(n798), .ip2(n786), .op(N899) );
  nor2_1 U1526 ( .ip1(n787), .ip2(n786), .op(N900) );
  nor2_1 U1527 ( .ip1(n788), .ip2(n786), .op(N901) );
  nor2_1 U1528 ( .ip1(n789), .ip2(n786), .op(N902) );
  nor2_1 U1529 ( .ip1(n790), .ip2(n786), .op(N903) );
  nor2_1 U1530 ( .ip1(n791), .ip2(n786), .op(N904) );
  nor2_1 U1531 ( .ip1(n792), .ip2(n786), .op(N905) );
  nor2_1 U1532 ( .ip1(n793), .ip2(n786), .op(N906) );
  nor2_1 U1533 ( .ip1(n794), .ip2(n786), .op(N907) );
  nor2_1 U1534 ( .ip1(n795), .ip2(n786), .op(N908) );
  nor2_1 U1535 ( .ip1(n800), .ip2(n786), .op(N909) );
  nor2_1 U1536 ( .ip1(n797), .ip2(n786), .op(N910) );
  nor2_1 U1537 ( .ip1(n781), .ip2(n786), .op(N911) );
  nand2_1 U1538 ( .ip1(w[12]), .ip2(n801), .op(n796) );
  nor2_1 U1539 ( .ip1(n798), .ip2(n796), .op(N915) );
  nor2_1 U1540 ( .ip1(n787), .ip2(n796), .op(N916) );
  nor2_1 U1541 ( .ip1(n788), .ip2(n796), .op(N917) );
  nor2_1 U1542 ( .ip1(n789), .ip2(n796), .op(N918) );
  nor2_1 U1543 ( .ip1(n790), .ip2(n796), .op(N919) );
  nor2_1 U1544 ( .ip1(n791), .ip2(n796), .op(N920) );
  nor2_1 U1545 ( .ip1(n792), .ip2(n796), .op(N921) );
  nor2_1 U1546 ( .ip1(n793), .ip2(n796), .op(N922) );
  nor2_1 U1547 ( .ip1(n794), .ip2(n796), .op(N923) );
  nor2_1 U1548 ( .ip1(n795), .ip2(n796), .op(N924) );
  nor2_1 U1549 ( .ip1(n800), .ip2(n796), .op(N925) );
  nor2_1 U1550 ( .ip1(n797), .ip2(n796), .op(N926) );
  nand2_1 U1551 ( .ip1(w[13]), .ip2(n801), .op(n799) );
  nor2_1 U1552 ( .ip1(n798), .ip2(n799), .op(N931) );
  nor2_1 U1553 ( .ip1(n787), .ip2(n799), .op(N932) );
  nor2_1 U1554 ( .ip1(n788), .ip2(n799), .op(N933) );
  nor2_1 U1555 ( .ip1(n789), .ip2(n799), .op(N934) );
  nor2_1 U1556 ( .ip1(n790), .ip2(n799), .op(N935) );
  nor2_1 U1557 ( .ip1(n791), .ip2(n799), .op(N936) );
  nor2_1 U1558 ( .ip1(n792), .ip2(n799), .op(N937) );
  nor2_1 U1559 ( .ip1(n793), .ip2(n799), .op(N938) );
  nor2_1 U1560 ( .ip1(n794), .ip2(n799), .op(N939) );
  nor2_1 U1561 ( .ip1(n795), .ip2(n799), .op(N940) );
  nor2_1 U1562 ( .ip1(n800), .ip2(n799), .op(N941) );
  nand2_1 U1563 ( .ip1(w[14]), .ip2(n801), .op(n802) );
  nor2_1 U1564 ( .ip1(n798), .ip2(n802), .op(N947) );
  nor2_1 U1565 ( .ip1(n787), .ip2(n802), .op(N948) );
  nor2_1 U1566 ( .ip1(n788), .ip2(n802), .op(N949) );
  nor2_1 U1567 ( .ip1(n789), .ip2(n802), .op(N950) );
  nor2_1 U1568 ( .ip1(n790), .ip2(n802), .op(N951) );
  nor2_1 U1569 ( .ip1(n791), .ip2(n802), .op(N952) );
  nor2_1 U1570 ( .ip1(n792), .ip2(n802), .op(N953) );
  nor2_1 U1571 ( .ip1(n793), .ip2(n802), .op(N954) );
  nor2_1 U1572 ( .ip1(n794), .ip2(n802), .op(N955) );
  nor2_1 U1573 ( .ip1(n795), .ip2(n802), .op(N956) );
  nor2_1 U1574 ( .ip1(\layer4[0][8] ), .ip2(\layer4[1][8] ), .op(n803) );
  nand2_1 U1575 ( .ip1(\layer4[0][8] ), .ip2(\layer4[1][8] ), .op(n804) );
  inv_1 U1576 ( .ip(n804), .op(n805) );
  nor3_1 U1577 ( .ip1(n803), .ip2(n483), .ip3(n805), .op(N707) );
  mux2_1 U1578 ( .ip1(n805), .ip2(n804), .s(\layer4[1][9] ), .op(n807) );
  nor2_1 U1579 ( .ip1(\layer4[0][9] ), .ip2(n807), .op(n806) );
  not_ab_or_c_or_d U1580 ( .ip1(\layer4[0][9] ), .ip2(n807), .ip3(reset), 
        .ip4(n806), .op(N708) );
  nand2_1 U1581 ( .ip1(\layer4[1][9] ), .ip2(\layer4[0][9] ), .op(n810) );
  or2_1 U1582 ( .ip1(\layer4[1][9] ), .ip2(\layer4[0][9] ), .op(n808) );
  nand3_1 U1583 ( .ip1(\layer4[1][8] ), .ip2(\layer4[0][8] ), .ip3(n808), .op(
        n809) );
  nand2_1 U1584 ( .ip1(n810), .ip2(n809), .op(n812) );
  and2_1 U1585 ( .ip1(n811), .ip2(n801), .op(N709) );
  fulladder U1586 ( .a(\layer4[1][10] ), .b(\layer4[0][10] ), .ci(n812), .co(
        n814), .s(n811) );
  and2_1 U1587 ( .ip1(n813), .ip2(n835), .op(N710) );
  fulladder U1588 ( .a(\layer4[1][11] ), .b(\layer4[0][11] ), .ci(n814), .co(
        n816), .s(n813) );
  and2_1 U1589 ( .ip1(n815), .ip2(n835), .op(N711) );
  fulladder U1590 ( .a(\layer4[1][12] ), .b(\layer4[0][12] ), .ci(n816), .co(
        n818), .s(n815) );
  and2_1 U1591 ( .ip1(n817), .ip2(n835), .op(N712) );
  fulladder U1592 ( .a(\layer4[1][13] ), .b(\layer4[0][13] ), .ci(n818), .co(
        n820), .s(n817) );
  and2_1 U1593 ( .ip1(n819), .ip2(n835), .op(N713) );
  fulladder U1594 ( .a(\layer4[1][14] ), .b(\layer4[0][14] ), .ci(n820), .co(
        n822), .s(n819) );
  and2_1 U1595 ( .ip1(n821), .ip2(n835), .op(N714) );
  fulladder U1596 ( .a(\layer4[1][15] ), .b(\layer4[0][15] ), .ci(n822), .co(
        n824), .s(n821) );
  and2_1 U1597 ( .ip1(n823), .ip2(n835), .op(N715) );
  fulladder U1598 ( .a(\layer4[1][16] ), .b(\layer4[0][16] ), .ci(n824), .co(
        n826), .s(n823) );
  and2_1 U1599 ( .ip1(n825), .ip2(n835), .op(N716) );
  fulladder U1600 ( .a(\layer4[1][17] ), .b(\layer4[0][17] ), .ci(n826), .co(
        n828), .s(n825) );
  and2_1 U1601 ( .ip1(n827), .ip2(n835), .op(N717) );
  fulladder U1602 ( .a(\layer4[1][18] ), .b(\layer4[0][18] ), .ci(n828), .co(
        n830), .s(n827) );
  and2_1 U1603 ( .ip1(n829), .ip2(n835), .op(N718) );
  fulladder U1604 ( .a(\layer4[1][19] ), .b(\layer4[0][19] ), .ci(n830), .co(
        n832), .s(n829) );
  and2_1 U1605 ( .ip1(n831), .ip2(n835), .op(N719) );
  fulladder U1606 ( .a(\layer4[1][20] ), .b(\layer4[0][20] ), .ci(n832), .co(
        n834), .s(n831) );
  and2_1 U1607 ( .ip1(n833), .ip2(n835), .op(N720) );
  fulladder U1608 ( .a(\layer4[1][21] ), .b(\layer4[0][21] ), .ci(n834), .co(
        n837), .s(n833) );
  and2_1 U1609 ( .ip1(n836), .ip2(n835), .op(N721) );
  fulladder U1610 ( .a(\layer4[1][22] ), .b(\layer4[0][22] ), .ci(n837), .co(
        n840), .s(n836) );
  xor2_1 U1611 ( .ip1(\layer4[1][23] ), .ip2(\layer4[0][23] ), .op(n839) );
  nor2_1 U1612 ( .ip1(n840), .ip2(n839), .op(n838) );
  not_ab_or_c_or_d U1613 ( .ip1(n840), .ip2(n839), .ip3(reset), .ip4(n838), 
        .op(N722) );
endmodule

